magic
tech sky130A
magscale 1 2
timestamp 1731213143
<< nwell >>
rect 5922 -1882 5926 -1832
rect 5596 -1884 5926 -1882
rect 5596 -1896 5828 -1884
rect 5596 -1898 5830 -1896
rect 5596 -1900 5920 -1898
rect 5922 -1900 5926 -1884
rect 5596 -2000 5926 -1900
<< locali >>
rect 5512 -1510 5650 -1502
rect 5512 -1544 5532 -1510
rect 5626 -1544 5650 -1510
rect 5512 -1562 5650 -1544
rect 5556 -1626 5604 -1562
rect 5954 -1784 6102 -1754
rect 5014 -1858 5082 -1848
rect 5014 -1968 5022 -1858
rect 5072 -1868 5082 -1858
rect 5118 -1868 5222 -1866
rect 5072 -1886 5222 -1868
rect 5556 -1886 5604 -1838
rect 5072 -1902 5292 -1886
rect 5392 -1902 5604 -1886
rect 5072 -1952 5604 -1902
rect 5698 -1884 5806 -1830
rect 5954 -1870 5988 -1784
rect 6066 -1854 6102 -1784
rect 6066 -1870 6104 -1854
rect 5698 -1896 5828 -1884
rect 5698 -1898 5830 -1896
rect 5698 -1900 5920 -1898
rect 5954 -1900 6104 -1870
rect 5698 -1944 6104 -1900
rect 5756 -1950 6104 -1944
rect 5072 -1954 5222 -1952
rect 5072 -1956 5128 -1954
rect 5072 -1968 5082 -1956
rect 5014 -1980 5082 -1968
rect 5928 -1962 6104 -1950
rect 5022 -2246 5372 -2234
rect 5022 -2382 5034 -2246
rect 5098 -2382 5372 -2246
rect 5928 -2292 6046 -1962
rect 5410 -2340 5702 -2296
rect 5774 -2340 6046 -2292
rect 5022 -2392 5372 -2382
rect 5282 -2944 5398 -2930
rect 5282 -3028 5288 -2944
rect 5396 -3028 5398 -2944
rect 5282 -3042 5398 -3028
rect 5898 -3110 6064 -3096
rect 5898 -3114 5918 -3110
rect 5486 -3160 5720 -3122
rect 5808 -3160 5918 -3114
rect 5898 -3188 5918 -3160
rect 6042 -3188 6064 -3110
rect 5898 -3200 6064 -3188
rect 5174 -3476 5590 -3444
rect 5174 -3518 5188 -3476
rect 5234 -3508 5590 -3476
rect 5234 -3518 5278 -3508
rect 5174 -3524 5278 -3518
rect 5376 -3524 5590 -3508
rect 5542 -3564 5590 -3524
rect 5542 -3836 5590 -3732
rect 5542 -3974 5592 -3836
rect 5536 -4176 5584 -4046
rect 5446 -4204 5702 -4176
rect 5446 -4288 5482 -4204
rect 5664 -4288 5702 -4204
rect 5446 -4312 5702 -4288
<< viali >>
rect 5532 -1544 5626 -1510
rect 5022 -1968 5072 -1858
rect 5988 -1870 6066 -1784
rect 5034 -2382 5098 -2246
rect 5288 -3028 5396 -2944
rect 5918 -3188 6042 -3110
rect 5188 -3518 5234 -3476
rect 5700 -3784 5748 -3746
rect 5482 -4288 5664 -4204
<< metal1 >>
rect 6090 -254 6322 -250
rect 5858 -260 6322 -254
rect 5858 -438 6090 -260
rect 6190 -438 6388 -260
rect 5858 -444 6388 -438
rect 5858 -450 6322 -444
rect 5858 -454 6160 -450
rect 5350 -564 6054 -558
rect 5350 -570 6196 -564
rect 5290 -582 6196 -570
rect 9858 -572 10132 -568
rect 9858 -574 10166 -572
rect 5290 -738 6136 -582
rect 6262 -738 6272 -582
rect 9660 -588 10166 -574
rect 5290 -752 6196 -738
rect 5290 -1402 5398 -752
rect 5854 -754 6098 -752
rect 5854 -758 6054 -754
rect 9660 -766 9758 -588
rect 9880 -766 10166 -588
rect 9660 -772 10166 -766
rect 9660 -788 10132 -772
rect 9660 -794 9934 -788
rect 5924 -802 6056 -798
rect 5924 -816 6440 -802
rect 5924 -900 5942 -816
rect 6040 -840 6440 -816
rect 6040 -900 6056 -840
rect 5924 -920 6056 -900
rect 5832 -1108 5934 -1106
rect 5832 -1150 6058 -1108
rect 5832 -1282 5960 -1150
rect 6046 -1282 6058 -1150
rect 5832 -1308 6058 -1282
rect 5280 -1598 5398 -1402
rect 5472 -1378 5672 -1328
rect 5832 -1332 5940 -1308
rect 5472 -1484 5522 -1378
rect 5640 -1484 5672 -1378
rect 5472 -1510 5672 -1484
rect 5472 -1528 5532 -1510
rect 5520 -1544 5532 -1528
rect 5626 -1528 5672 -1510
rect 5838 -1494 5940 -1332
rect 5626 -1544 5638 -1528
rect 5520 -1556 5638 -1544
rect 5838 -1592 5936 -1494
rect 5142 -1800 5220 -1796
rect 4974 -1846 5106 -1806
rect 4974 -1986 5014 -1846
rect 5086 -1986 5106 -1846
rect 4974 -2010 5106 -1986
rect 5142 -1862 5320 -1800
rect 4986 -2246 5114 -2212
rect 4986 -2272 5034 -2246
rect 5098 -2272 5114 -2246
rect 4986 -2362 4998 -2272
rect 5106 -2362 5114 -2272
rect 4986 -2382 5034 -2362
rect 5098 -2382 5114 -2362
rect 4986 -2416 5114 -2382
rect 5142 -2508 5220 -1862
rect 5520 -2060 5614 -1964
rect 5836 -1970 5930 -1832
rect 5962 -1898 5968 -1758
rect 6110 -1898 6120 -1758
rect 5836 -2062 6068 -1970
rect 5912 -2064 6068 -2062
rect 5140 -2602 5282 -2508
rect 5140 -2604 5230 -2602
rect 5504 -2604 5634 -2506
rect 5140 -2636 5226 -2604
rect 5140 -2892 5246 -2636
rect 5548 -2882 5632 -2784
rect 5928 -2786 6066 -2064
rect 5888 -2878 6294 -2786
rect 5140 -3072 5238 -2892
rect 5270 -2932 5416 -2926
rect 5270 -2944 5428 -2932
rect 5270 -2946 5288 -2944
rect 5396 -2946 5428 -2944
rect 5266 -3030 5276 -2946
rect 5418 -3030 5428 -2946
rect 5270 -3040 5428 -3030
rect 6186 -3040 6294 -2878
rect 5270 -3046 5416 -3040
rect 6182 -3064 6294 -3040
rect 5140 -3322 5246 -3072
rect 5890 -3108 6078 -3088
rect 5890 -3186 5916 -3108
rect 5890 -3188 5918 -3186
rect 6042 -3188 6078 -3108
rect 5890 -3206 6078 -3188
rect 5140 -3404 5316 -3322
rect 5140 -3422 5372 -3404
rect 5146 -3426 5372 -3422
rect 5552 -3424 5634 -3326
rect 5552 -3426 5598 -3424
rect 5146 -3432 5246 -3426
rect 5180 -3474 5250 -3464
rect 5128 -3476 5250 -3474
rect 5128 -3480 5188 -3476
rect 5234 -3480 5250 -3476
rect 5122 -3600 5132 -3480
rect 5244 -3514 5254 -3480
rect 5244 -3600 5250 -3514
rect 5282 -3570 5372 -3426
rect 5626 -3458 5790 -3452
rect 5626 -3552 5636 -3458
rect 5784 -3552 5794 -3458
rect 5902 -3546 6148 -3542
rect 6182 -3546 6290 -3064
rect 5626 -3558 5790 -3552
rect 5126 -3608 5250 -3600
rect 5684 -3654 5752 -3558
rect 5902 -3630 6292 -3546
rect 6046 -3634 6292 -3630
rect 5682 -3686 5752 -3654
rect 5680 -3702 5752 -3686
rect 5680 -3740 5750 -3702
rect 5680 -3746 5760 -3740
rect 5680 -3764 5700 -3746
rect 5686 -3784 5700 -3764
rect 5748 -3784 5760 -3746
rect 5686 -3788 5760 -3784
rect 5686 -3800 5756 -3788
rect 5276 -3870 5374 -3806
rect 5820 -3874 5916 -3808
rect 5456 -4192 5694 -4180
rect 5456 -4296 5466 -4192
rect 5682 -4296 5694 -4192
rect 5456 -4306 5694 -4296
<< via1 >>
rect 6090 -438 6190 -260
rect 6136 -738 6262 -582
rect 9758 -766 9880 -588
rect 5942 -900 6040 -816
rect 5960 -1282 6046 -1150
rect 5522 -1484 5640 -1378
rect 5014 -1858 5086 -1846
rect 5014 -1968 5022 -1858
rect 5022 -1968 5072 -1858
rect 5072 -1968 5086 -1858
rect 5014 -1986 5086 -1968
rect 4998 -2362 5034 -2272
rect 5034 -2362 5098 -2272
rect 5098 -2362 5106 -2272
rect 5968 -1784 6110 -1758
rect 5968 -1870 5988 -1784
rect 5988 -1870 6066 -1784
rect 6066 -1870 6110 -1784
rect 5968 -1898 6110 -1870
rect 5276 -3028 5288 -2946
rect 5288 -3028 5396 -2946
rect 5396 -3028 5418 -2946
rect 5276 -3030 5418 -3028
rect 5916 -3110 6042 -3108
rect 5916 -3186 5918 -3110
rect 5918 -3186 6042 -3110
rect 5132 -3518 5188 -3480
rect 5188 -3518 5234 -3480
rect 5234 -3518 5244 -3480
rect 5132 -3600 5244 -3518
rect 5636 -3552 5784 -3458
rect 5466 -4204 5682 -4192
rect 5466 -4288 5482 -4204
rect 5482 -4288 5664 -4204
rect 5664 -4288 5682 -4204
rect 5466 -4296 5682 -4288
<< metal2 >>
rect 9992 252 10156 268
rect 9992 174 10014 252
rect 9994 148 10014 174
rect 10130 174 10156 252
rect 10130 148 10154 174
rect 9994 114 10154 148
rect 6090 -260 6190 -250
rect 6190 -276 6294 -266
rect 9486 -296 9734 -240
rect 9486 -324 9554 -296
rect 6190 -438 6294 -430
rect 6090 -440 6294 -438
rect 7124 -406 9554 -324
rect 9686 -406 9734 -296
rect 6090 -448 6190 -440
rect 7124 -468 9734 -406
rect 7124 -478 9586 -468
rect 6138 -562 6294 -552
rect 6136 -582 6138 -572
rect 6136 -748 6138 -738
rect 6138 -762 6294 -752
rect 7124 -754 7256 -478
rect 9660 -588 9934 -574
rect 7122 -786 7270 -754
rect 5924 -816 6056 -798
rect 5924 -900 5942 -816
rect 6040 -900 6056 -816
rect 5924 -920 6056 -900
rect 7124 -1022 7270 -786
rect 9660 -766 9758 -588
rect 9882 -766 9934 -588
rect 9660 -794 9934 -766
rect 7122 -1134 7270 -1022
rect 5950 -1138 6316 -1136
rect 6720 -1138 7270 -1134
rect 5950 -1150 7270 -1138
rect 5950 -1286 5960 -1150
rect 6046 -1152 7270 -1150
rect 6046 -1272 6188 -1152
rect 6338 -1266 7270 -1152
rect 6338 -1272 6470 -1266
rect 6046 -1286 6470 -1272
rect 6656 -1286 7270 -1266
rect 5950 -1296 6316 -1286
rect 7122 -1288 7270 -1286
rect 9664 -904 9824 -900
rect 9994 -904 10152 114
rect 9664 -1142 10156 -904
rect 5490 -1378 5654 -1366
rect 5490 -1492 5506 -1378
rect 5640 -1484 5654 -1378
rect 5636 -1492 5654 -1484
rect 5490 -1508 5654 -1492
rect 5960 -1480 6110 -1460
rect 5960 -1594 5982 -1480
rect 6078 -1594 6110 -1480
rect 5960 -1758 6110 -1594
rect 5960 -1776 5968 -1758
rect 5014 -1846 5086 -1836
rect 5086 -1980 5248 -1848
rect 5968 -1908 6110 -1898
rect 5086 -1986 5236 -1980
rect 5014 -1988 5236 -1986
rect 5014 -1996 5086 -1988
rect 5128 -2018 5236 -1988
rect 4998 -2272 5106 -2262
rect 4998 -2372 5106 -2362
rect 5000 -3468 5106 -2372
rect 5138 -2948 5236 -2018
rect 5952 -2374 7210 -2370
rect 9664 -2374 9824 -1142
rect 9994 -1146 10152 -1142
rect 5942 -2376 7210 -2374
rect 9370 -2376 9824 -2374
rect 5942 -2462 9824 -2376
rect 5942 -2470 7200 -2462
rect 9370 -2464 9824 -2462
rect 5942 -2894 6026 -2470
rect 5928 -2920 6026 -2894
rect 5276 -2946 5418 -2936
rect 5138 -3030 5276 -2948
rect 5138 -3032 5418 -3030
rect 5138 -3036 5236 -3032
rect 5276 -3040 5418 -3032
rect 5928 -3098 6014 -2920
rect 5916 -3108 6042 -3098
rect 5914 -3186 5916 -3174
rect 5914 -3188 6042 -3186
rect 5912 -3438 6042 -3188
rect 5634 -3458 6042 -3438
rect 5000 -3470 5138 -3468
rect 5000 -3480 5244 -3470
rect 5000 -3600 5132 -3480
rect 5634 -3552 5636 -3458
rect 5784 -3504 6042 -3458
rect 5924 -3508 6042 -3504
rect 5634 -3556 5784 -3552
rect 5636 -3562 5784 -3556
rect 5000 -3610 5244 -3600
rect 5000 -3614 5138 -3610
rect 5096 -3616 5138 -3614
rect 5456 -4192 5694 -4180
rect 5456 -4296 5466 -4192
rect 5682 -4296 5694 -4192
rect 5456 -4306 5694 -4296
<< via2 >>
rect 10014 148 10130 252
rect 6102 -430 6190 -276
rect 6190 -430 6294 -276
rect 9554 -406 9686 -296
rect 6138 -582 6294 -562
rect 6138 -738 6262 -582
rect 6262 -738 6294 -582
rect 6138 -752 6294 -738
rect 5942 -900 6040 -816
rect 9760 -766 9880 -588
rect 9880 -766 9882 -588
rect 5960 -1282 6046 -1154
rect 6188 -1272 6338 -1152
rect 5960 -1286 6046 -1282
rect 5506 -1484 5522 -1378
rect 5522 -1484 5636 -1378
rect 5506 -1492 5636 -1484
rect 5982 -1594 6078 -1480
rect 5466 -4296 5682 -4192
<< metal3 >>
rect 8022 1330 8838 1462
rect 8588 14 8786 1330
rect 10004 252 10140 257
rect 8916 238 9114 252
rect 10004 250 10014 252
rect 9578 240 10014 250
rect 8862 216 9114 238
rect 9476 216 10014 240
rect 8862 148 10014 216
rect 10130 148 10140 252
rect 8862 146 10140 148
rect 8862 142 9518 146
rect 10004 143 10140 146
rect 8588 -86 8744 14
rect 6062 -242 6330 -230
rect 6062 -258 6574 -242
rect 8588 -258 8734 -86
rect 8862 -170 8922 142
rect 6062 -262 8734 -258
rect 6062 -276 8744 -262
rect 6062 -430 6102 -276
rect 6294 -292 8744 -276
rect 6294 -298 8752 -292
rect 6294 -300 8788 -298
rect 8930 -300 9088 -258
rect 6294 -302 9088 -300
rect 6294 -430 6790 -302
rect 6062 -444 6790 -430
rect 6954 -312 9088 -302
rect 6954 -444 8868 -312
rect 6062 -464 8868 -444
rect 9068 -464 9088 -312
rect 6062 -466 9088 -464
rect 6306 -478 9088 -466
rect 9486 -292 9734 -240
rect 9486 -406 9554 -292
rect 9686 -406 9734 -292
rect 9486 -468 9734 -406
rect 6538 -546 9436 -544
rect 6118 -562 9436 -546
rect 6118 -752 6138 -562
rect 6294 -582 9436 -562
rect 6294 -600 9202 -582
rect 6294 -732 6478 -600
rect 6640 -712 9202 -600
rect 6640 -718 6904 -712
rect 6640 -732 6768 -718
rect 6294 -752 6768 -732
rect 7112 -740 9202 -712
rect 6118 -768 6768 -752
rect 6432 -772 6768 -768
rect 7122 -752 9202 -740
rect 9384 -752 9436 -582
rect 7122 -772 9436 -752
rect 9660 -588 9934 -574
rect 9660 -602 9760 -588
rect 7122 -774 7380 -772
rect 7122 -786 7276 -774
rect 5926 -800 6030 -798
rect 5926 -816 6060 -800
rect 5926 -900 5942 -816
rect 6040 -900 6060 -816
rect 5926 -920 6060 -900
rect 5978 -950 6060 -920
rect 5978 -992 6062 -950
rect 5772 -1000 6062 -992
rect 5768 -1044 6062 -1000
rect 7124 -1022 7276 -786
rect 9660 -780 9688 -602
rect 9882 -766 9934 -588
rect 9810 -780 9934 -766
rect 9660 -794 9934 -780
rect 9660 -804 9922 -794
rect 7110 -1034 7276 -1022
rect 5768 -1056 6060 -1044
rect 5768 -1070 5856 -1056
rect 5458 -1378 5692 -1322
rect 5458 -1492 5506 -1378
rect 5636 -1492 5692 -1378
rect 5768 -1384 5854 -1070
rect 5968 -1149 6090 -1126
rect 5950 -1154 6090 -1149
rect 5950 -1286 5960 -1154
rect 6046 -1286 6090 -1154
rect 5950 -1291 6090 -1286
rect 5968 -1312 6090 -1291
rect 6168 -1152 6366 -1138
rect 6168 -1282 6188 -1152
rect 6338 -1272 6366 -1152
rect 6320 -1282 6366 -1272
rect 6168 -1304 6366 -1282
rect 5768 -1448 6090 -1384
rect 5770 -1480 6090 -1448
rect 5770 -1486 5982 -1480
rect 5458 -4080 5692 -1492
rect 5968 -1574 5982 -1486
rect 5972 -1594 5982 -1574
rect 6078 -1574 6090 -1480
rect 6078 -1594 6088 -1574
rect 5972 -1599 6088 -1594
rect 7050 -1666 7276 -1034
rect 7064 -1962 7276 -1666
rect 7050 -2356 7276 -1962
rect 7014 -2366 7522 -2356
rect 7014 -2368 7558 -2366
rect 7656 -2368 7766 -2364
rect 7014 -2478 7766 -2368
rect 7050 -2484 7766 -2478
rect 7050 -2488 7558 -2484
rect 7656 -2500 7766 -2484
rect 5456 -4086 5692 -4080
rect 5456 -4160 5690 -4086
rect 5450 -4192 5696 -4160
rect 5450 -4296 5466 -4192
rect 5682 -4296 5696 -4192
rect 5450 -4310 5696 -4296
<< via3 >>
rect 6790 -444 6954 -302
rect 8868 -464 9068 -312
rect 9554 -296 9686 -292
rect 9554 -406 9686 -296
rect 6478 -732 6640 -600
rect 9202 -752 9384 -582
rect 9688 -766 9760 -602
rect 9760 -766 9810 -602
rect 9688 -780 9810 -766
rect 6188 -1272 6320 -1172
rect 6188 -1282 6320 -1272
<< metal4 >>
rect 9734 -186 9735 -180
rect 6752 -302 6990 -258
rect 6752 -444 6790 -302
rect 6954 -444 6990 -302
rect 6440 -600 6678 -546
rect 6440 -732 6478 -600
rect 6640 -732 6678 -600
rect 6440 -792 6678 -732
rect 6752 -816 6990 -444
rect 7836 -812 8006 -218
rect 8850 -312 9086 -222
rect 9176 -232 9416 -190
rect 8850 -464 8868 -312
rect 9068 -464 9086 -312
rect 8850 -482 9086 -464
rect 9174 -582 9416 -232
rect 9484 -292 9734 -194
rect 9484 -406 9554 -292
rect 9686 -406 9734 -292
rect 9484 -422 9734 -406
rect 9486 -468 9734 -422
rect 9174 -752 9202 -582
rect 9384 -734 9416 -582
rect 9672 -602 9840 -576
rect 9384 -752 9414 -734
rect 9174 -776 9414 -752
rect 9672 -780 9688 -602
rect 9810 -780 9840 -602
rect 6187 -1172 6321 -1171
rect 6187 -1282 6188 -1172
rect 6320 -1282 6321 -1172
rect 9672 -1184 9840 -780
rect 6187 -1283 6321 -1282
rect 7944 -1358 9840 -1184
rect 9672 -1368 9840 -1358
use tt_asw_3v3  x1
timestamp 1731213143
transform 1 0 6104 0 1 -5137
box 0 -757 10957 4352
use tt_asw_3v3  x2
timestamp 1731213143
transform -1 0 9755 0 -1 4116
box 0 -757 10957 4352
use sky130_fd_sc_hd__inv_1  x3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5536 0 1 -2556
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  x4 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 0 1 5340 1 0 -1864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1704896540
transform 0 1 5320 1 0 -4138
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  x6
timestamp 1704896540
transform 0 1 5326 1 0 -3818
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1704896540
transform -1 0 5880 0 1 -2556
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x8
timestamp 1704896540
transform -1 0 5568 0 1 -3378
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1704896540
transform -1 0 5900 0 1 -3376
box -38 -48 314 592
<< labels >>
flabel metal1 5858 -454 6058 -254 0 FreeSans 256 0 0 0 VDDA
port 1 nsew
flabel metal1 5854 -758 6054 -558 0 FreeSans 256 0 0 0 GND
port 0 nsew
flabel metal1 9966 -772 10166 -572 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
flabel metal1 5858 -1308 6058 -1108 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 5472 -1528 5672 -1328 0 FreeSans 256 0 0 0 Cin
port 2 nsew
<< end >>
