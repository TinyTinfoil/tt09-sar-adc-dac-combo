magic
tech sky130A
magscale 1 2
timestamp 1731252669
<< metal1 >>
rect 20543 44763 20745 44769
rect 20543 43893 20745 44561
rect 10913 43691 20745 43893
rect 822 38628 1178 38698
rect 822 38364 832 38628
rect 1134 38616 1178 38628
rect 1804 38616 2020 38617
rect 1134 38402 3206 38616
rect 8016 38574 8584 38587
rect 1134 38364 1178 38402
rect 822 38332 1178 38364
rect 786 34580 1236 34736
rect 786 34318 874 34580
rect 1100 34576 1236 34580
rect 1804 34576 2020 38402
rect 8016 38372 9118 38574
rect 8348 38360 9118 38372
rect 8568 37206 8976 38360
rect 8568 36870 8614 37206
rect 8910 36870 8976 37206
rect 8568 36794 8976 36870
rect 1100 34318 2054 34576
rect 786 34293 2054 34318
rect 786 34194 1236 34293
rect 1804 28668 2020 34293
rect 8058 28668 8508 28675
rect 1804 28452 3318 28668
rect 8058 28460 9128 28668
rect 8358 28454 9128 28460
rect 1806 23080 2018 28452
rect 8578 27300 8986 28454
rect 8578 26964 8624 27300
rect 8920 26964 8986 27300
rect 8578 26888 8986 26964
rect 798 22910 1242 23066
rect 798 22648 880 22910
rect 1106 22906 1242 22910
rect 1806 22906 2026 23080
rect 1106 22648 2050 22906
rect 798 22623 2050 22648
rect 798 22524 1242 22623
rect 1806 22520 2026 22623
rect 1806 20690 2018 22520
rect 1806 20394 2030 20690
rect 1806 19036 2018 20394
rect 1806 18824 3422 19036
rect 8314 19030 8522 19036
rect 1809 13834 2016 18824
rect 8314 18816 9228 19030
rect 8314 18814 8522 18816
rect 8678 17662 9086 18816
rect 8678 17326 8724 17662
rect 9020 17326 9086 17662
rect 8678 17250 9086 17326
rect 4123 14069 4325 14075
rect 10913 14069 11115 43691
rect 26608 38587 27047 44611
rect 20118 38582 20500 38586
rect 19500 38384 20500 38582
rect 25400 38405 27047 38587
rect 19500 38368 20270 38384
rect 19642 37214 20050 38368
rect 19642 36878 19708 37214
rect 20004 36878 20050 37214
rect 19642 36802 20050 36878
rect 26608 28685 27047 38405
rect 20034 28660 20590 28670
rect 19474 28468 20590 28660
rect 25328 28491 27047 28685
rect 19474 28446 20244 28468
rect 19616 27292 20024 28446
rect 19616 26956 19682 27292
rect 19978 26956 20024 27292
rect 19616 26880 20024 26956
rect 26608 18905 27047 28491
rect 19994 18872 20634 18878
rect 19492 18676 20634 18872
rect 25328 18711 27047 18905
rect 19492 18658 20262 18676
rect 19634 17504 20042 18658
rect 19634 17168 19700 17504
rect 19996 17168 20042 17504
rect 19634 17092 20042 17168
rect 4325 13867 11115 14069
rect 4123 13861 4325 13867
rect 1806 13538 2022 13834
rect 1809 12674 2016 13538
rect 792 12504 1236 12660
rect 792 12242 874 12504
rect 1100 12500 1236 12504
rect 1804 12500 2020 12674
rect 1100 12242 2044 12500
rect 792 12217 2044 12242
rect 792 12118 1236 12217
rect 1804 12114 2020 12217
rect 1809 8971 2016 12114
rect 1766 8922 2058 8971
rect 1766 8715 3373 8922
rect 1766 2671 2058 8715
rect 8188 8696 9126 8910
rect 19876 8906 20450 8938
rect 26608 8925 27047 18711
rect 8576 7542 8984 8696
rect 19290 8692 20450 8906
rect 25196 8731 27047 8925
rect 8576 7206 8622 7542
rect 8918 7206 8984 7542
rect 8576 7130 8984 7206
rect 19432 7538 19840 8692
rect 19876 8682 20450 8692
rect 19432 7202 19498 7538
rect 19794 7202 19840 7538
rect 19432 7126 19840 7202
rect 26608 2671 27047 8731
rect 1698 2242 27047 2671
rect 26608 2237 27047 2242
<< via1 >>
rect 20543 44561 20745 44763
rect 832 38364 1134 38628
rect 874 34318 1100 34580
rect 8614 36870 8910 37206
rect 8624 26964 8920 27300
rect 880 22648 1106 22910
rect 8724 17326 9020 17662
rect 19708 36878 20004 37214
rect 19682 26956 19978 27292
rect 19700 17168 19996 17504
rect 4123 13867 4325 14069
rect 874 12242 1100 12504
rect 8622 7206 8918 7542
rect 19498 7202 19794 7538
<< metal2 >>
rect 20543 44891 20745 44900
rect 15090 44575 15099 44777
rect 15301 44575 15310 44777
rect 21679 44811 21881 44820
rect 11379 44136 11388 44371
rect 11623 44136 11632 44371
rect 832 38628 1134 38638
rect 832 38354 1134 38364
rect 220 38078 568 38112
rect 220 37858 252 38078
rect 526 38052 568 38078
rect 526 38044 1232 38052
rect 526 37858 3424 38044
rect 220 37852 3424 37858
rect 220 37810 568 37852
rect 1034 37848 3424 37852
rect 826 34580 1156 34628
rect 826 34318 874 34580
rect 1100 34318 1156 34580
rect 826 34270 1156 34318
rect 204 30794 596 30836
rect 204 30572 242 30794
rect 544 30753 596 30794
rect 1997 30753 2187 37848
rect 8532 37262 9140 37288
rect 8486 37252 9186 37262
rect 8486 36594 9186 36604
rect 11388 36051 11623 44136
rect 12234 43729 12243 43931
rect 12445 43729 12454 43931
rect 7947 35816 11623 36051
rect 7947 33691 8182 35816
rect 12243 34997 12445 43729
rect 10775 34795 12445 34997
rect 7944 33469 7953 33691
rect 8175 33469 8184 33691
rect 7947 33463 8182 33469
rect 544 30572 2187 30753
rect 204 30563 2187 30572
rect 204 30546 596 30563
rect 1997 28155 2187 30563
rect 1997 27965 3481 28155
rect 832 22910 1162 22958
rect 832 22648 880 22910
rect 1106 22648 1162 22910
rect 832 22600 1162 22648
rect 2000 20690 2184 27965
rect 8542 27356 9150 27382
rect 8496 27346 9196 27356
rect 8496 26688 9196 26698
rect 3023 23937 3215 23941
rect 10775 23937 10977 34795
rect 3018 23932 10977 23937
rect 3018 23740 3023 23932
rect 3215 23740 10977 23932
rect 3018 23735 10977 23740
rect 3023 23731 3215 23735
rect 15099 21903 15301 44575
rect 20537 44561 20543 44763
rect 20745 44561 20751 44763
rect 21679 43759 21881 44609
rect 23347 44225 23549 44234
rect 25950 44225 26142 44229
rect 23549 44220 26147 44225
rect 23549 44028 25950 44220
rect 26142 44028 26147 44220
rect 23549 44023 26147 44028
rect 23347 44014 23549 44023
rect 25950 44019 26142 44023
rect 20107 43557 21881 43759
rect 23941 43869 24143 43878
rect 25531 43869 25723 43873
rect 24143 43864 25728 43869
rect 24143 43672 25531 43864
rect 25723 43672 25728 43864
rect 24143 43667 25728 43672
rect 23941 43658 24143 43667
rect 25531 43663 25723 43667
rect 20107 40991 20309 43557
rect 16621 40789 20309 40991
rect 16621 23877 16823 40789
rect 26463 38037 26961 44627
rect 25130 37853 26961 38037
rect 19478 37270 20086 37296
rect 19432 37260 20132 37270
rect 19432 36602 20132 36612
rect 26463 28123 26961 37853
rect 25158 27939 26961 28123
rect 19452 27348 20060 27374
rect 19406 27338 20106 27348
rect 19406 26680 20106 26690
rect 24752 23877 24944 23881
rect 16621 23872 24949 23877
rect 16621 23680 24752 23872
rect 24944 23680 24949 23872
rect 16621 23675 24949 23680
rect 24752 23671 24944 23675
rect 15099 21701 16713 21903
rect 214 20642 606 20684
rect 214 20420 252 20642
rect 554 20601 606 20642
rect 2000 20601 2197 20690
rect 554 20420 2197 20601
rect 214 20411 2197 20420
rect 214 20394 606 20411
rect 2000 20394 2197 20411
rect 2000 18486 2184 20394
rect 2000 18302 3614 18486
rect 2003 13834 2182 18302
rect 8642 17718 9250 17744
rect 8596 17708 9296 17718
rect 8596 17050 9296 17060
rect 2952 14064 4123 14069
rect 2948 13872 2957 14064
rect 3149 13872 4123 14064
rect 2952 13867 4123 13872
rect 4325 13867 4331 14069
rect 16511 14047 16713 21701
rect 26463 18343 26961 27939
rect 25154 18159 26961 18343
rect 19470 17560 20078 17586
rect 19424 17550 20124 17560
rect 19424 16892 20124 16902
rect 25399 14047 25591 14051
rect 16511 14042 25596 14047
rect 16511 13850 25399 14042
rect 25591 13850 25596 14042
rect 16511 13845 25596 13850
rect 25399 13841 25591 13845
rect 206 13786 598 13828
rect 206 13564 244 13786
rect 546 13745 598 13786
rect 1999 13745 2189 13834
rect 546 13564 2189 13745
rect 206 13555 2189 13564
rect 206 13538 598 13555
rect 1999 13538 2189 13555
rect 826 12504 1156 12552
rect 826 12242 874 12504
rect 1100 12242 1156 12504
rect 826 12194 1156 12242
rect 2003 8431 2182 13538
rect 1968 8396 2217 8431
rect 1968 8217 3517 8396
rect 26463 8363 26961 18159
rect 1968 2778 2217 8217
rect 25002 8179 26961 8363
rect 8540 7598 9148 7624
rect 8494 7588 9194 7598
rect 19268 7594 19876 7620
rect 8494 6930 9194 6940
rect 19222 7584 19922 7594
rect 19222 6926 19922 6936
rect 26463 2778 26961 8179
rect 1844 2282 26961 2778
rect 26463 2281 26961 2282
<< via2 >>
rect 15099 44575 15301 44777
rect 20543 44763 20745 44891
rect 11388 44136 11623 44371
rect 832 38364 1134 38628
rect 252 37858 526 38078
rect 874 34318 1100 34580
rect 242 30572 544 30794
rect 8486 37206 9186 37252
rect 8486 36870 8614 37206
rect 8614 36870 8910 37206
rect 8910 36870 9186 37206
rect 8486 36604 9186 36870
rect 12243 43729 12445 43931
rect 7953 33469 8175 33691
rect 880 22648 1106 22910
rect 8496 27300 9196 27346
rect 8496 26964 8624 27300
rect 8624 26964 8920 27300
rect 8920 26964 9196 27300
rect 8496 26698 9196 26964
rect 3023 23740 3215 23932
rect 20543 44689 20745 44763
rect 21679 44609 21881 44811
rect 23347 44023 23549 44225
rect 25950 44028 26142 44220
rect 23941 43667 24143 43869
rect 25531 43672 25723 43864
rect 19432 37214 20132 37260
rect 19432 36878 19708 37214
rect 19708 36878 20004 37214
rect 20004 36878 20132 37214
rect 19432 36612 20132 36878
rect 19406 27292 20106 27338
rect 19406 26956 19682 27292
rect 19682 26956 19978 27292
rect 19978 26956 20106 27292
rect 19406 26690 20106 26956
rect 24752 23680 24944 23872
rect 252 20420 554 20642
rect 8596 17662 9296 17708
rect 8596 17326 8724 17662
rect 8724 17326 9020 17662
rect 9020 17326 9296 17662
rect 8596 17060 9296 17326
rect 2957 13872 3149 14064
rect 19424 17504 20124 17550
rect 19424 17168 19700 17504
rect 19700 17168 19996 17504
rect 19996 17168 20124 17504
rect 19424 16902 20124 17168
rect 25399 13850 25591 14042
rect 244 13564 546 13786
rect 874 12242 1100 12504
rect 8494 7542 9194 7588
rect 8494 7206 8622 7542
rect 8622 7206 8918 7542
rect 8918 7206 9194 7542
rect 8494 6940 9194 7206
rect 19222 7538 19922 7584
rect 19222 7202 19498 7538
rect 19498 7202 19794 7538
rect 19794 7202 19922 7538
rect 19222 6936 19922 7202
<< metal3 >>
rect 20543 45009 20745 45015
rect 15094 44777 15306 44782
rect 15094 44575 15099 44777
rect 15301 44575 15655 44777
rect 15857 44575 15863 44777
rect 20538 44689 20543 44896
rect 21679 44931 21881 44937
rect 20745 44689 20750 44896
rect 20538 44684 20750 44689
rect 21674 44609 21679 44816
rect 22278 44828 22448 44886
rect 21881 44609 21886 44816
rect 22278 44646 22320 44828
rect 21674 44604 21886 44609
rect 15094 44570 15306 44575
rect 22252 44512 22320 44646
rect 22414 44646 22448 44828
rect 22798 44826 22968 44884
rect 22798 44689 22840 44826
rect 22414 44545 22460 44646
rect 22414 44512 22499 44545
rect 11383 44371 11628 44376
rect 22252 44371 22499 44512
rect 11383 44136 11388 44371
rect 11623 44136 22499 44371
rect 22771 44510 22840 44689
rect 22934 44689 22968 44826
rect 23360 44814 23530 44872
rect 22934 44662 22973 44689
rect 23360 44668 23402 44814
rect 22934 44510 22986 44662
rect 22771 44264 22986 44510
rect 23352 44498 23402 44668
rect 23496 44668 23530 44814
rect 23926 44798 24088 44842
rect 23496 44498 23560 44668
rect 23352 44430 23560 44498
rect 23926 44472 23962 44798
rect 24058 44472 24088 44798
rect 23352 44413 23580 44430
rect 11383 44131 11628 44136
rect 12238 43931 12450 43936
rect 22771 43931 22973 44264
rect 23347 44230 23580 44413
rect 23926 44349 24088 44472
rect 24476 44790 24640 44826
rect 24476 44440 24500 44790
rect 24608 44440 24640 44790
rect 23926 44328 24143 44349
rect 23342 44228 23580 44230
rect 23342 44225 23554 44228
rect 23342 44023 23347 44225
rect 23549 44023 23554 44225
rect 23342 44018 23554 44023
rect 23924 44010 24143 44328
rect 12238 43729 12243 43931
rect 12445 43729 22973 43931
rect 23898 43874 24143 44010
rect 23898 43869 24148 43874
rect 12238 43724 12450 43729
rect 23898 43667 23941 43869
rect 24143 43667 24148 43869
rect 23898 43662 24148 43667
rect 23898 43624 24026 43662
rect 2864 43512 3042 43514
rect 24476 43512 24640 44440
rect 25945 44220 26741 44225
rect 25945 44028 25950 44220
rect 26142 44028 26741 44220
rect 25945 44023 26741 44028
rect 25526 43864 25728 43883
rect 25526 43672 25531 43864
rect 25723 43672 25728 43864
rect 2864 43304 24662 43512
rect 822 38628 1144 38633
rect 822 38364 832 38628
rect 1134 38364 1144 38628
rect 822 38359 1144 38364
rect 242 38078 536 38083
rect 242 37858 252 38078
rect 526 37858 536 38078
rect 242 37853 536 37858
rect 2864 37630 3042 43304
rect 16862 39900 18240 40724
rect 19064 39900 19070 40724
rect 8348 37266 10548 39466
rect 18070 37274 20270 39474
rect 25526 37637 25728 43672
rect 8448 37252 9248 37266
rect 8448 36604 8486 37252
rect 9186 36604 9248 37252
rect 19370 37260 20170 37274
rect 8448 36466 9248 36604
rect 10532 35968 11426 36792
rect 12250 35968 12256 36792
rect 19370 36612 19432 37260
rect 20132 36612 20170 37260
rect 19370 36474 20170 36612
rect 10532 35206 11356 35968
rect 826 34580 1156 34628
rect 826 34318 874 34580
rect 1100 34318 1156 34580
rect 826 34270 1156 34318
rect 26539 34129 26741 44023
rect 25526 33927 26741 34129
rect 2296 33691 8318 33696
rect 2296 33469 7953 33691
rect 8175 33469 8318 33691
rect 2296 33464 8318 33469
rect 232 30794 554 30799
rect 232 30572 242 30794
rect 544 30572 554 30794
rect 232 30567 554 30572
rect 2296 27925 2528 33464
rect 16854 30220 20242 31028
rect 2296 27723 3088 27925
rect 2296 27708 2528 27723
rect 8358 27360 10558 29560
rect 16854 28422 17662 30220
rect 16854 27608 17662 27614
rect 8458 27346 9258 27360
rect 18044 27352 20244 29552
rect 25526 27723 25728 33927
rect 8458 26698 8496 27346
rect 9196 26698 9258 27346
rect 8458 26560 9258 26698
rect 19344 27338 20144 27352
rect 19344 26690 19406 27338
rect 20106 26690 20144 27338
rect 19344 26552 20144 26690
rect 10442 26350 11250 26356
rect 10442 25536 11250 25542
rect 3018 23932 3220 23937
rect 3018 23740 3023 23932
rect 3215 23740 3220 23932
rect 832 22910 1162 22958
rect 832 22648 880 22910
rect 1106 22648 1162 22910
rect 832 22600 1162 22648
rect 242 20642 564 20647
rect 242 20420 252 20642
rect 554 20420 564 20642
rect 242 20415 564 20420
rect 3018 18077 3220 23740
rect 24747 23872 25728 23877
rect 24747 23680 24752 23872
rect 24944 23680 25728 23872
rect 24747 23675 25728 23680
rect 16692 21018 17516 21024
rect 17516 20194 20160 21018
rect 16692 20188 17516 20194
rect 8458 17722 10658 19922
rect 8558 17708 9358 17722
rect 8558 17060 8596 17708
rect 9296 17060 9358 17708
rect 18062 17564 20262 19764
rect 25526 17943 25728 23675
rect 8558 16922 9358 17060
rect 19362 17550 20162 17564
rect 19362 16902 19424 17550
rect 20124 16902 20162 17550
rect 19362 16764 20162 16902
rect 8454 15554 9262 15560
rect 2952 14064 3154 14069
rect 2952 13872 2957 14064
rect 3149 13872 3154 14064
rect 234 13786 556 13791
rect 234 13564 244 13786
rect 546 13564 556 13786
rect 234 13559 556 13564
rect 826 12504 1156 12552
rect 826 12242 874 12504
rect 1100 12242 1156 12504
rect 826 12194 1156 12242
rect 2952 7963 3154 13872
rect 8454 10518 9262 14746
rect 19266 12338 20074 14274
rect 25394 14042 25596 14047
rect 25394 13850 25399 14042
rect 25591 13850 25596 14042
rect 19260 11530 19266 12338
rect 20074 11530 20080 12338
rect 17860 7598 20060 9798
rect 25394 7963 25596 13850
rect 8484 7588 9204 7593
rect 8484 6940 8494 7588
rect 9194 6940 9204 7588
rect 8484 6935 9204 6940
rect 19160 7584 19960 7598
rect 19160 6936 19222 7584
rect 19922 6936 19960 7584
rect 19160 6798 19960 6936
rect 9536 3690 9546 4420
rect 10204 3690 10214 4420
rect 17990 4309 18930 4310
rect 17955 3371 17961 4309
rect 18959 3371 18965 4309
rect 17990 1606 18930 3371
rect 17990 1394 27350 1606
rect 17990 964 26720 1394
rect 27150 964 27350 1394
rect 17990 666 27350 964
<< via3 >>
rect 15655 44575 15857 44777
rect 20543 44891 20745 45009
rect 20543 44807 20745 44891
rect 21679 44811 21881 44931
rect 21679 44729 21881 44811
rect 22320 44512 22414 44828
rect 22840 44510 22934 44826
rect 23402 44498 23496 44814
rect 23962 44472 24058 44798
rect 24500 44440 24608 44790
rect 832 38364 1134 38628
rect 252 37858 526 38078
rect 18240 39900 19064 40724
rect 11426 35968 12250 36792
rect 874 34318 1100 34580
rect 242 30572 544 30794
rect 16854 27614 17662 28422
rect 10442 25542 11250 26350
rect 880 22648 1106 22910
rect 252 20420 554 20642
rect 16692 20194 17516 21018
rect 8454 14746 9262 15554
rect 244 13564 546 13786
rect 874 12242 1100 12504
rect 19266 11530 20074 12338
rect 9546 3690 10204 4420
rect 17961 3371 18959 4309
rect 26720 964 27150 1394
<< mimcap >>
rect 8448 38366 10448 39366
rect 8448 37466 9548 38366
rect 10348 37466 10448 38366
rect 8448 37366 10448 37466
rect 18170 38374 20170 39374
rect 18170 37474 18270 38374
rect 19070 37474 20170 38374
rect 18170 37374 20170 37474
rect 8458 28460 10458 29460
rect 8458 27560 9558 28460
rect 10358 27560 10458 28460
rect 8458 27460 10458 27560
rect 18144 28452 20144 29452
rect 18144 27552 18244 28452
rect 19044 27552 20144 28452
rect 18144 27452 20144 27552
rect 8558 18822 10558 19822
rect 8558 17922 9658 18822
rect 10458 17922 10558 18822
rect 8558 17822 10558 17922
rect 18162 18664 20162 19664
rect 18162 17764 18262 18664
rect 19062 17764 20162 18664
rect 18162 17664 20162 17764
rect 17960 8698 19960 9698
rect 17960 7798 18060 8698
rect 18860 7798 19960 8698
rect 17960 7698 19960 7798
<< mimcapcontact >>
rect 9548 37466 10348 38366
rect 18270 37474 19070 38374
rect 9558 27560 10358 28460
rect 18244 27552 19044 28452
rect 9658 17922 10458 18822
rect 18262 17764 19062 18664
rect 18060 7798 18860 8698
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20543 45010 20745 45157
rect 21222 45109 21282 45152
rect 20542 45009 20746 45010
rect 20542 44807 20543 45009
rect 20745 44807 20746 45009
rect 20542 44806 20746 44807
rect 15654 44777 15858 44778
rect 15654 44575 15655 44777
rect 15857 44575 20017 44777
rect 15654 44574 15858 44575
rect 200 38078 600 44152
rect 200 37858 252 38078
rect 526 37858 600 38078
rect 200 30794 600 37858
rect 200 30572 242 30794
rect 544 30572 600 30794
rect 200 20690 600 30572
rect 800 38628 1200 44152
rect 800 38364 832 38628
rect 1134 38364 1200 38628
rect 800 34580 1200 38364
rect 800 34318 874 34580
rect 1100 34318 1200 34580
rect 800 23080 1200 34318
rect 1400 38880 1800 44152
rect 19815 44097 20017 44575
rect 21105 44097 21307 45109
rect 21679 44932 21881 45169
rect 22326 45010 22386 45152
rect 22878 45010 22938 45152
rect 21678 44931 21882 44932
rect 21678 44729 21679 44931
rect 21881 44729 21882 44931
rect 22282 44828 22442 45010
rect 22282 44808 22320 44828
rect 21678 44728 21882 44729
rect 22284 44512 22320 44808
rect 22414 44512 22442 44828
rect 22284 44466 22442 44512
rect 22804 44848 22958 45010
rect 23430 44996 23490 45152
rect 23982 45038 24042 45152
rect 22804 44826 22962 44848
rect 23368 44836 23522 44996
rect 22804 44510 22840 44826
rect 22934 44510 22962 44826
rect 22804 44464 22962 44510
rect 23366 44814 23524 44836
rect 23366 44498 23402 44814
rect 23496 44498 23524 44814
rect 23366 44452 23524 44498
rect 23926 44798 24086 45038
rect 24534 45012 24594 45152
rect 23926 44472 23962 44798
rect 24058 44472 24086 44798
rect 23926 44344 24086 44472
rect 24476 44790 24642 45012
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 24476 44440 24500 44790
rect 24608 44440 24642 44790
rect 24476 44336 24642 44440
rect 19815 43895 21307 44097
rect 9528 40916 12708 41916
rect 1400 38714 3732 38880
rect 1400 28970 1800 38714
rect 9528 38466 10528 40916
rect 18239 40724 19065 40725
rect 18239 39900 18240 40724
rect 19064 39900 19065 40724
rect 18239 39899 19065 39900
rect 18240 38474 19064 39899
rect 26373 38875 26784 44643
rect 24838 38707 26784 38875
rect 9448 38366 10528 38466
rect 9448 37466 9548 38366
rect 10348 37802 10528 38366
rect 18170 38374 19170 38474
rect 10348 37466 10448 37802
rect 9448 37278 10448 37466
rect 18170 37474 18270 38374
rect 19070 37474 19170 38374
rect 9436 36793 11708 37278
rect 9436 36792 12251 36793
rect 9436 36454 11426 36792
rect 10884 35968 11426 36454
rect 12250 35968 12251 36792
rect 18170 36474 19170 37474
rect 11425 35967 12251 35968
rect 18242 35434 19063 36474
rect 1400 28798 3770 28970
rect 1400 23080 1800 28798
rect 9340 28560 10340 31056
rect 26373 28961 26784 38707
rect 24814 28793 26784 28961
rect 9340 28460 10458 28560
rect 9340 27560 9558 28460
rect 10358 27560 10458 28460
rect 18144 28452 19144 28552
rect 16853 28422 17663 28423
rect 18144 28422 18244 28452
rect 16853 27614 16854 28422
rect 17662 27614 18244 28422
rect 16853 27613 17663 27614
rect 9340 27402 10458 27560
rect 18144 27552 18244 27614
rect 19044 27552 19144 28452
rect 9340 27400 11250 27402
rect 9458 26560 11250 27400
rect 10442 26351 11250 26560
rect 10441 26350 11251 26351
rect 10441 25542 10442 26350
rect 11250 25542 11251 26350
rect 10441 25541 11251 25542
rect 18144 25300 19144 27552
rect 800 22910 1206 23080
rect 800 22648 880 22910
rect 1106 22648 1206 22910
rect 800 22520 1206 22648
rect 1400 22520 1806 23080
rect 800 20690 1200 22520
rect 1400 20690 1800 22520
rect 200 20642 610 20690
rect 200 20420 252 20642
rect 554 20420 610 20642
rect 200 20394 610 20420
rect 800 20394 1210 20690
rect 1400 20394 1810 20690
rect 200 13834 600 20394
rect 800 13834 1200 20394
rect 1400 19302 1800 20394
rect 1396 19130 3766 19302
rect 1400 13834 1800 19130
rect 9554 18922 10342 21206
rect 16691 21018 17517 21019
rect 16691 20194 16692 21018
rect 17516 20194 17517 21018
rect 16691 20193 17517 20194
rect 16692 19504 17516 20193
rect 9554 18822 10558 18922
rect 9554 18468 9658 18822
rect 9558 17922 9658 18468
rect 10458 17922 10558 18822
rect 16692 18680 19204 19504
rect 26373 19181 26784 28793
rect 24838 19013 26784 19181
rect 9558 16922 10558 17922
rect 18162 18664 19204 18680
rect 18162 17764 18262 18664
rect 19062 17828 19204 18664
rect 19062 17764 19162 17828
rect 8453 15554 9263 15555
rect 9746 15554 10554 16922
rect 8453 14746 8454 15554
rect 9262 14746 10554 15554
rect 8453 14745 9263 14746
rect 18162 14490 19162 17764
rect 200 13786 602 13834
rect 200 13564 244 13786
rect 546 13564 602 13786
rect 200 13538 602 13564
rect 800 13538 1202 13834
rect 1400 13538 1802 13834
rect 200 1000 600 13538
rect 800 12504 1200 13538
rect 800 12242 874 12504
rect 1100 12242 1200 12504
rect 800 1000 1200 12242
rect 1400 9208 1800 13538
rect 1400 9036 3776 9208
rect 1400 2790 1800 9036
rect 9416 7960 10426 12550
rect 19265 12338 20075 12339
rect 18026 11530 19266 12338
rect 20074 11530 20075 12338
rect 18026 8798 18834 11530
rect 19265 11529 20075 11530
rect 26373 9201 26784 19013
rect 24650 9033 26784 9201
rect 17960 8698 18960 8798
rect 17960 7798 18060 8698
rect 18860 7798 18960 8698
rect 9514 7078 10290 7098
rect 8222 2790 9258 5328
rect 9478 4420 10290 7078
rect 9478 3690 9546 4420
rect 10204 3690 10290 4420
rect 9478 3664 10290 3690
rect 17960 4309 18960 7798
rect 9478 3644 10254 3664
rect 17960 3371 17961 4309
rect 18959 3371 18960 4309
rect 17960 3370 18960 3371
rect 26373 2790 26784 9033
rect 1400 2388 26784 2790
rect 1400 1000 1800 2388
rect 8222 2266 9258 2388
rect 26373 2384 26784 2388
rect 26478 1394 27406 1602
rect 26478 964 26720 1394
rect 27150 964 27406 1394
rect 26478 200 27406 964
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 26478 138 27414 200
rect 27234 0 27414 138
use dacswitch  dacswitch_0
timestamp 1731231864
transform 1 0 -1940 0 1 39157
box 4430 -5137 10166 4116
use dacswitch  dacswitch_1
timestamp 1731231864
transform -1 0 30554 0 1 39157
box 4430 -5137 10166 4116
use dacswitch  dacswitch_2
timestamp 1731231864
transform 1 0 -1940 0 1 29243
box 4430 -5137 10166 4116
use dacswitch  dacswitch_3
timestamp 1731231864
transform -1 0 30554 0 1 29243
box 4430 -5137 10166 4116
use dacswitch  dacswitch_4
timestamp 1731231864
transform 1 0 -1808 0 1 19597
box 4430 -5137 10166 4116
use dacswitch  dacswitch_5
timestamp 1731231864
transform -1 0 30554 0 1 19463
box 4430 -5137 10166 4116
use dacswitch  dacswitch_6
timestamp 1731231864
transform 1 0 -1874 0 1 9483
box 4430 -5137 10166 4116
use dacswitch  dacswitch_7
timestamp 1731231864
transform -1 0 30422 0 1 9483
box 4430 -5137 10166 4116
use mim400  mim400_0
timestamp 1731238228
transform 1 0 18142 0 1 30204
box -736 0 2216 5982
use mim400  mim400_1
timestamp 1731238228
transform 1 0 9150 0 -1 26366
box -736 0 2216 5982
use mim400  mim400_2
timestamp 1731238228
transform 1 0 9240 0 1 30056
box -736 0 2216 5982
use mim400  mim400_3
timestamp 1731238228
transform 0 -1 20266 -1 0 15566
box -736 0 2216 5982
use mim400  mim400_4
timestamp 1731238228
transform 1 0 18044 0 -1 26172
box -736 0 2216 5982
use mim400  mim400_5
timestamp 1731238228
transform 0 1 8438 -1 0 12618
box -736 0 2216 5982
use mim400  mim400_6
timestamp 1731238228
transform 0 1 11708 -1 0 42016
box -736 0 2216 5982
use mimcaptut200b  mimcaptut200b_0
timestamp 1731226444
transform -1 0 8456 0 1 8502
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_1
timestamp 1731226444
transform 1 0 10298 0 1 5258
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_2
timestamp 1731226444
transform -1 0 8558 0 1 18622
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_3
timestamp 1731226444
transform -1 0 8458 0 1 28260
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_4
timestamp 1731226444
transform -1 0 8448 0 1 38166
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_5
timestamp 1731226444
transform 1 0 19960 0 1 8498
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_6
timestamp 1731226444
transform 1 0 20170 0 1 38174
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_7
timestamp 1731226444
transform 1 0 20144 0 1 28252
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_8
timestamp 1731226444
transform 1 0 20162 0 1 18464
box -2100 -1700 100 1300
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
rlabel metal4 10058 16922 10058 16922 5 top
rlabel metal3 8958 16922 8958 16922 5 bot
rlabel metal4 9958 26560 9958 26560 5 top
rlabel metal3 8858 26560 8858 26560 5 bot
rlabel metal4 9948 36466 9948 36466 5 top
rlabel metal3 8848 36466 8848 36466 5 bot
rlabel metal4 18670 36474 18670 36474 5 top
rlabel metal3 19770 36474 19770 36474 5 bot
rlabel metal4 18644 26552 18644 26552 5 top
rlabel metal3 19744 26552 19744 26552 5 bot
rlabel metal4 18662 16764 18662 16764 5 top
rlabel metal3 19762 16764 19762 16764 5 bot
rlabel metal4 18460 6798 18460 6798 5 top
rlabel metal3 19560 6798 19560 6798 5 bot
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
