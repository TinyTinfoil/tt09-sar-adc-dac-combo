magic
tech sky130A
magscale 1 2
timestamp 1731231864
<< nwell >>
rect 5604 -1882 5608 -1832
rect 5278 -1884 5608 -1882
rect 5278 -1896 5510 -1884
rect 4432 -2000 4602 -1896
rect 5278 -1898 5512 -1896
rect 5278 -1900 5602 -1898
rect 5604 -1900 5608 -1884
rect 5278 -2000 5608 -1900
rect 4432 -2246 4960 -2000
rect 5216 -2218 5268 -2092
rect 4432 -2360 4602 -2246
rect 4430 -2820 4600 -2644
rect 4430 -2898 4988 -2820
rect 4430 -3056 5012 -2898
rect 4430 -3108 4600 -3056
rect 5262 -4154 5398 -4080
rect 5488 -4154 5596 -4136
rect 5262 -4204 5596 -4154
rect 5262 -4376 5598 -4204
rect 5040 -4534 5598 -4376
rect 5040 -4544 5592 -4534
rect 5040 -4546 5504 -4544
<< nsubdiff >>
rect 4471 -1967 4508 -1933
rect 4471 -1993 4505 -1967
rect 4471 -2289 4505 -2263
rect 4471 -2323 4508 -2289
rect 4469 -2715 4506 -2681
rect 4469 -2741 4503 -2715
rect 4469 -3037 4503 -3011
rect 4469 -3071 4506 -3037
rect 5432 -4415 5498 -4414
rect 5077 -4449 5137 -4415
rect 5407 -4449 5498 -4415
rect 5077 -4452 5111 -4449
rect 5432 -4450 5498 -4449
rect 5433 -4452 5467 -4450
<< nsubdiffcont >>
rect 4471 -2263 4505 -1993
rect 4469 -3011 4503 -2741
rect 5137 -4449 5407 -4415
<< locali >>
rect 5194 -1510 5332 -1502
rect 5194 -1544 5214 -1510
rect 5308 -1544 5332 -1510
rect 5194 -1562 5332 -1544
rect 5238 -1626 5286 -1562
rect 5636 -1784 5784 -1754
rect 4696 -1858 4764 -1848
rect 4471 -1967 4508 -1933
rect 4471 -1993 4505 -1967
rect 4696 -1968 4704 -1858
rect 4754 -1868 4764 -1858
rect 4800 -1868 4904 -1866
rect 4754 -1886 4904 -1868
rect 5238 -1886 5286 -1838
rect 4754 -1902 4974 -1886
rect 5074 -1902 5286 -1886
rect 4754 -1952 5286 -1902
rect 5380 -1884 5488 -1830
rect 5636 -1870 5670 -1784
rect 5748 -1854 5784 -1784
rect 5748 -1870 5786 -1854
rect 5380 -1896 5510 -1884
rect 5380 -1898 5512 -1896
rect 5380 -1900 5602 -1898
rect 5636 -1900 5786 -1870
rect 5380 -1944 5786 -1900
rect 5438 -1950 5786 -1944
rect 4754 -1954 4904 -1952
rect 4754 -1956 4810 -1954
rect 4754 -1968 4764 -1956
rect 4696 -1980 4764 -1968
rect 5610 -1962 5786 -1950
rect 4468 -2263 4471 -2182
rect 4816 -2070 4920 -2064
rect 4505 -2094 4920 -2070
rect 4505 -2172 4832 -2094
rect 4894 -2172 4920 -2094
rect 4505 -2188 4920 -2172
rect 4505 -2190 4890 -2188
rect 4505 -2263 4510 -2190
rect 4468 -2741 4510 -2263
rect 4704 -2246 5054 -2234
rect 4704 -2382 4716 -2246
rect 4780 -2382 5054 -2246
rect 5610 -2292 5728 -1962
rect 5092 -2340 5384 -2296
rect 5456 -2340 5728 -2292
rect 4704 -2392 5054 -2382
rect 4468 -2832 4469 -2741
rect 4503 -2832 4510 -2741
rect 4469 -3037 4503 -3011
rect 4964 -2944 5080 -2930
rect 4964 -3028 4970 -2944
rect 5078 -3028 5080 -2944
rect 4469 -3071 4506 -3037
rect 4964 -3042 5080 -3028
rect 5580 -3110 5746 -3096
rect 5580 -3114 5600 -3110
rect 5168 -3160 5402 -3122
rect 5490 -3160 5600 -3114
rect 5580 -3188 5600 -3160
rect 5724 -3188 5746 -3110
rect 5580 -3200 5746 -3188
rect 4856 -3476 5272 -3444
rect 4856 -3518 4870 -3476
rect 4916 -3508 5272 -3476
rect 4916 -3518 4960 -3508
rect 4856 -3524 4960 -3518
rect 5058 -3524 5272 -3508
rect 5224 -3564 5272 -3524
rect 5224 -3836 5272 -3732
rect 5224 -3974 5274 -3836
rect 4982 -4416 5018 -4076
rect 5218 -4176 5266 -4046
rect 5128 -4204 5384 -4176
rect 5128 -4288 5164 -4204
rect 5346 -4288 5384 -4204
rect 5128 -4312 5384 -4288
rect 5432 -4415 5498 -4414
rect 5077 -4416 5137 -4415
rect 4982 -4449 5137 -4416
rect 5407 -4449 5498 -4415
rect 4982 -4452 5111 -4449
rect 5432 -4450 5498 -4449
rect 5433 -4452 5467 -4450
rect 4982 -4458 5108 -4452
rect 4984 -4460 5108 -4458
<< viali >>
rect 5214 -1544 5308 -1510
rect 4704 -1968 4754 -1858
rect 5670 -1870 5748 -1784
rect 4832 -2172 4894 -2094
rect 4716 -2382 4780 -2246
rect 4970 -3028 5078 -2944
rect 5600 -3188 5724 -3110
rect 4870 -3518 4916 -3476
rect 5382 -3784 5430 -3746
rect 5164 -4288 5346 -4204
<< metal1 >>
rect 6090 -254 6322 -250
rect 5858 -260 6322 -254
rect 5858 -438 6090 -260
rect 6190 -438 6388 -260
rect 5858 -444 6388 -438
rect 5858 -450 6322 -444
rect 5858 -454 6160 -450
rect 5736 -558 6180 -554
rect 5032 -570 6180 -558
rect 4972 -588 6180 -570
rect 9858 -572 10132 -568
rect 9858 -574 10166 -572
rect 4972 -714 5988 -588
rect 6114 -714 6180 -588
rect 4972 -752 6180 -714
rect 4972 -1402 5080 -752
rect 5536 -756 6180 -752
rect 9660 -588 10166 -574
rect 5536 -758 5736 -756
rect 9660 -766 9758 -588
rect 9880 -766 10166 -588
rect 9660 -772 10166 -766
rect 9660 -788 10132 -772
rect 9660 -794 9934 -788
rect 5606 -802 5738 -798
rect 5778 -802 6162 -798
rect 5606 -816 6440 -802
rect 5606 -900 5624 -816
rect 5722 -840 6440 -816
rect 5722 -900 5738 -840
rect 5778 -842 6162 -840
rect 5606 -920 5738 -900
rect 5514 -1108 5616 -1106
rect 5514 -1150 5740 -1108
rect 5514 -1282 5642 -1150
rect 5728 -1282 5740 -1150
rect 5514 -1308 5740 -1282
rect 4962 -1598 5080 -1402
rect 5154 -1378 5354 -1328
rect 5514 -1332 5622 -1308
rect 5154 -1484 5204 -1378
rect 5322 -1484 5354 -1378
rect 5154 -1510 5354 -1484
rect 5154 -1528 5214 -1510
rect 5202 -1544 5214 -1528
rect 5308 -1528 5354 -1510
rect 5520 -1494 5622 -1332
rect 5308 -1544 5320 -1528
rect 5202 -1556 5320 -1544
rect 5520 -1592 5618 -1494
rect 4824 -1800 4902 -1796
rect 4656 -1846 4788 -1806
rect 4656 -1986 4696 -1846
rect 4768 -1986 4788 -1846
rect 4656 -2010 4788 -1986
rect 4824 -1862 5002 -1800
rect 4824 -2094 4902 -1862
rect 5202 -2060 5296 -1964
rect 5518 -1970 5612 -1832
rect 5644 -1898 5650 -1758
rect 5792 -1898 5802 -1758
rect 5518 -2062 5750 -1970
rect 5594 -2064 5750 -2062
rect 4824 -2172 4832 -2094
rect 4894 -2172 4902 -2094
rect 4668 -2246 4796 -2212
rect 4668 -2272 4716 -2246
rect 4780 -2272 4796 -2246
rect 4668 -2362 4680 -2272
rect 4788 -2362 4796 -2272
rect 4668 -2382 4716 -2362
rect 4780 -2382 4796 -2362
rect 4668 -2416 4796 -2382
rect 4824 -2508 4902 -2172
rect 4822 -2602 4964 -2508
rect 4822 -2604 4912 -2602
rect 5186 -2604 5316 -2506
rect 4822 -2636 4908 -2604
rect 4822 -2892 4928 -2636
rect 5610 -2756 5748 -2064
rect 5610 -2784 5778 -2756
rect 5230 -2882 5314 -2784
rect 5610 -2786 6204 -2784
rect 5570 -2878 6294 -2786
rect 4822 -3072 4920 -2892
rect 4952 -2932 5098 -2926
rect 4952 -2944 5110 -2932
rect 4952 -2946 4970 -2944
rect 5078 -2946 5110 -2944
rect 4948 -3030 4958 -2946
rect 5100 -3030 5110 -2946
rect 4952 -3040 5110 -3030
rect 6186 -3040 6294 -2878
rect 4952 -3046 5098 -3040
rect 6182 -3064 6294 -3040
rect 4822 -3322 4928 -3072
rect 5572 -3108 5760 -3088
rect 5572 -3186 5598 -3108
rect 5572 -3188 5600 -3186
rect 5724 -3188 5760 -3108
rect 5572 -3206 5760 -3188
rect 4822 -3404 4998 -3322
rect 4822 -3422 5054 -3404
rect 4828 -3426 5054 -3422
rect 5234 -3424 5316 -3326
rect 5234 -3426 5280 -3424
rect 4828 -3432 4928 -3426
rect 4862 -3474 4932 -3464
rect 4810 -3476 4932 -3474
rect 4810 -3480 4870 -3476
rect 4916 -3480 4932 -3476
rect 4804 -3600 4814 -3480
rect 4926 -3514 4936 -3480
rect 4926 -3600 4932 -3514
rect 4964 -3570 5054 -3426
rect 5308 -3458 5472 -3452
rect 5308 -3552 5318 -3458
rect 5466 -3552 5476 -3458
rect 6182 -3536 6290 -3064
rect 5920 -3540 6290 -3536
rect 5812 -3542 6290 -3540
rect 5584 -3546 6290 -3542
rect 5308 -3558 5472 -3552
rect 4808 -3608 4932 -3600
rect 5366 -3654 5434 -3558
rect 5584 -3630 6292 -3546
rect 5728 -3634 6292 -3630
rect 5812 -3636 6156 -3634
rect 5364 -3686 5434 -3654
rect 5362 -3702 5434 -3686
rect 5362 -3740 5432 -3702
rect 5362 -3746 5442 -3740
rect 5362 -3764 5382 -3746
rect 5368 -3784 5382 -3764
rect 5430 -3784 5442 -3746
rect 5368 -3788 5442 -3784
rect 5368 -3800 5438 -3788
rect 4958 -3870 5056 -3806
rect 5502 -3874 5598 -3808
rect 5138 -4192 5376 -4180
rect 5138 -4296 5148 -4192
rect 5364 -4296 5376 -4192
rect 5138 -4306 5376 -4296
<< via1 >>
rect 6090 -438 6190 -260
rect 5988 -714 6114 -588
rect 9758 -766 9880 -588
rect 5624 -900 5722 -816
rect 5642 -1282 5728 -1150
rect 5204 -1484 5322 -1378
rect 4696 -1858 4768 -1846
rect 4696 -1968 4704 -1858
rect 4704 -1968 4754 -1858
rect 4754 -1968 4768 -1858
rect 4696 -1986 4768 -1968
rect 5650 -1784 5792 -1758
rect 5650 -1870 5670 -1784
rect 5670 -1870 5748 -1784
rect 5748 -1870 5792 -1784
rect 5650 -1898 5792 -1870
rect 4680 -2362 4716 -2272
rect 4716 -2362 4780 -2272
rect 4780 -2362 4788 -2272
rect 4958 -3028 4970 -2946
rect 4970 -3028 5078 -2946
rect 5078 -3028 5100 -2946
rect 4958 -3030 5100 -3028
rect 5598 -3110 5724 -3108
rect 5598 -3186 5600 -3110
rect 5600 -3186 5724 -3110
rect 4814 -3518 4870 -3480
rect 4870 -3518 4916 -3480
rect 4916 -3518 4926 -3480
rect 4814 -3600 4926 -3518
rect 5318 -3552 5466 -3458
rect 5148 -4204 5364 -4192
rect 5148 -4288 5164 -4204
rect 5164 -4288 5346 -4204
rect 5346 -4288 5364 -4204
rect 5148 -4296 5364 -4288
<< metal2 >>
rect 9992 252 10156 268
rect 9992 174 10014 252
rect 9994 148 10014 174
rect 10130 174 10156 252
rect 10130 148 10154 174
rect 9994 114 10154 148
rect 6090 -260 6190 -250
rect 6190 -276 6294 -266
rect 9486 -296 9734 -240
rect 9486 -324 9554 -296
rect 6190 -438 6294 -430
rect 6090 -440 6294 -438
rect 7124 -406 9554 -324
rect 9686 -406 9734 -296
rect 6090 -448 6190 -440
rect 7124 -468 9734 -406
rect 7124 -478 9586 -468
rect 5988 -584 6114 -578
rect 5984 -588 6114 -584
rect 5984 -594 5988 -588
rect 6110 -720 6114 -714
rect 5984 -724 6114 -720
rect 5984 -730 6110 -724
rect 7124 -754 7256 -478
rect 9660 -588 9934 -574
rect 7122 -786 7270 -754
rect 5606 -816 5738 -798
rect 5606 -900 5624 -816
rect 5722 -900 5738 -816
rect 5606 -920 5738 -900
rect 7124 -1022 7270 -786
rect 9660 -766 9758 -588
rect 9882 -766 9934 -588
rect 9660 -794 9934 -766
rect 5212 -1128 5572 -1120
rect 5212 -1136 5670 -1128
rect 5800 -1136 6172 -1132
rect 7122 -1134 7270 -1022
rect 5212 -1138 6316 -1136
rect 6720 -1138 7270 -1134
rect 5212 -1150 7270 -1138
rect 5212 -1286 5642 -1150
rect 5728 -1152 7270 -1150
rect 5728 -1272 6188 -1152
rect 6338 -1266 7270 -1152
rect 6338 -1272 6470 -1266
rect 5728 -1286 6470 -1272
rect 6656 -1286 7270 -1266
rect 5212 -1292 6316 -1286
rect 7122 -1288 7270 -1286
rect 9664 -904 9824 -900
rect 9994 -904 10152 114
rect 9664 -1142 10156 -904
rect 5212 -1296 5824 -1292
rect 6142 -1296 6316 -1292
rect 5212 -1302 5670 -1296
rect 5212 -1304 5572 -1302
rect 5172 -1378 5336 -1366
rect 5172 -1492 5188 -1378
rect 5322 -1484 5336 -1378
rect 5318 -1492 5336 -1484
rect 5172 -1508 5336 -1492
rect 5642 -1480 5792 -1460
rect 5642 -1594 5664 -1480
rect 5760 -1594 5792 -1480
rect 5642 -1758 5792 -1594
rect 5642 -1776 5650 -1758
rect 4696 -1846 4768 -1836
rect 4768 -1980 4930 -1848
rect 5650 -1908 5792 -1898
rect 4768 -1986 4918 -1980
rect 4696 -1988 4918 -1986
rect 4696 -1996 4768 -1988
rect 4810 -2018 4918 -1988
rect 4680 -2272 4788 -2262
rect 4680 -2372 4788 -2362
rect 4682 -3468 4788 -2372
rect 4820 -2948 4918 -2018
rect 5788 -2370 6168 -2368
rect 5634 -2374 7210 -2370
rect 9664 -2374 9824 -1142
rect 9994 -1146 10152 -1142
rect 5624 -2376 7210 -2374
rect 9370 -2376 9824 -2374
rect 5624 -2462 9824 -2376
rect 5624 -2470 7200 -2462
rect 9370 -2464 9824 -2462
rect 5624 -2894 5708 -2470
rect 5788 -2472 6168 -2470
rect 5610 -2920 5708 -2894
rect 4958 -2946 5100 -2936
rect 4820 -3030 4958 -2948
rect 4820 -3032 5100 -3030
rect 4820 -3036 4918 -3032
rect 4958 -3040 5100 -3032
rect 5610 -3098 5696 -2920
rect 5598 -3108 5724 -3098
rect 5596 -3186 5598 -3174
rect 5596 -3188 5724 -3186
rect 5594 -3438 5724 -3188
rect 5316 -3458 5724 -3438
rect 4682 -3470 4820 -3468
rect 4682 -3480 4926 -3470
rect 4682 -3600 4814 -3480
rect 5316 -3552 5318 -3458
rect 5466 -3504 5724 -3458
rect 5606 -3508 5724 -3504
rect 5316 -3556 5466 -3552
rect 5318 -3562 5466 -3556
rect 4682 -3610 4926 -3600
rect 4682 -3614 4820 -3610
rect 4778 -3616 4820 -3614
rect 5138 -4192 5376 -4180
rect 5138 -4296 5148 -4192
rect 5364 -4296 5376 -4192
rect 5138 -4306 5376 -4296
<< via2 >>
rect 10014 148 10130 252
rect 6102 -430 6190 -276
rect 6190 -430 6294 -276
rect 9554 -406 9686 -296
rect 5984 -714 5988 -594
rect 5988 -714 6110 -594
rect 5984 -720 6110 -714
rect 5624 -900 5722 -816
rect 9760 -766 9880 -588
rect 9880 -766 9882 -588
rect 5642 -1282 5728 -1154
rect 6188 -1272 6338 -1152
rect 5642 -1286 5728 -1282
rect 5188 -1484 5204 -1378
rect 5204 -1484 5318 -1378
rect 5188 -1492 5318 -1484
rect 5664 -1594 5760 -1480
rect 5148 -4296 5364 -4192
<< metal3 >>
rect 8022 1330 8838 1462
rect 8588 14 8786 1330
rect 10004 252 10140 257
rect 8916 238 9114 252
rect 10004 250 10014 252
rect 9578 240 10014 250
rect 8862 216 9114 238
rect 9476 216 10014 240
rect 8862 148 10014 216
rect 10130 148 10140 252
rect 8862 146 10140 148
rect 8862 142 9518 146
rect 10004 143 10140 146
rect 8588 -86 8744 14
rect 6062 -242 6330 -230
rect 6062 -258 6574 -242
rect 8588 -258 8734 -86
rect 8862 -170 8922 142
rect 6062 -262 8734 -258
rect 6062 -276 8744 -262
rect 6062 -430 6102 -276
rect 6294 -292 8744 -276
rect 6294 -298 8752 -292
rect 6294 -300 8788 -298
rect 8930 -300 9088 -258
rect 6294 -302 9088 -300
rect 6294 -430 6790 -302
rect 6062 -444 6790 -430
rect 6954 -312 9088 -302
rect 6954 -444 8868 -312
rect 6062 -464 8868 -444
rect 9068 -464 9088 -312
rect 6062 -466 9088 -464
rect 6306 -478 9088 -466
rect 9486 -292 9734 -240
rect 9486 -406 9554 -292
rect 9686 -406 9734 -292
rect 9486 -468 9734 -406
rect 6538 -546 9436 -544
rect 5974 -582 9436 -546
rect 5974 -594 9202 -582
rect 5974 -720 5984 -594
rect 6110 -600 9202 -594
rect 6110 -720 6478 -600
rect 5974 -732 6478 -720
rect 6640 -712 9202 -600
rect 6640 -718 6904 -712
rect 6640 -732 6768 -718
rect 5974 -762 6768 -732
rect 7112 -740 9202 -712
rect 6322 -768 6768 -762
rect 6432 -772 6768 -768
rect 7122 -752 9202 -740
rect 9384 -752 9436 -582
rect 7122 -772 9436 -752
rect 9660 -588 9934 -574
rect 9660 -602 9760 -588
rect 7122 -774 7380 -772
rect 7122 -786 7276 -774
rect 5608 -800 5712 -798
rect 5608 -816 5742 -800
rect 5608 -900 5624 -816
rect 5722 -900 5742 -816
rect 5608 -920 5742 -900
rect 5660 -950 5742 -920
rect 5660 -992 5744 -950
rect 5454 -1000 5744 -992
rect 5450 -1044 5744 -1000
rect 7124 -1022 7276 -786
rect 9660 -780 9688 -602
rect 9882 -766 9934 -588
rect 9810 -780 9934 -766
rect 9660 -794 9934 -780
rect 9660 -804 9922 -794
rect 7110 -1034 7276 -1022
rect 5450 -1056 5742 -1044
rect 5450 -1070 5538 -1056
rect 4826 -1322 5372 -1318
rect 4826 -1378 5374 -1322
rect 4826 -1492 5188 -1378
rect 5318 -1492 5374 -1378
rect 5450 -1384 5536 -1070
rect 5650 -1149 5772 -1126
rect 5632 -1154 5772 -1149
rect 5632 -1286 5642 -1154
rect 5728 -1286 5772 -1154
rect 5632 -1291 5772 -1286
rect 5650 -1312 5772 -1291
rect 6168 -1152 6366 -1138
rect 6168 -1282 6188 -1152
rect 6338 -1272 6366 -1152
rect 6320 -1282 6366 -1272
rect 6168 -1304 6366 -1282
rect 5450 -1448 5772 -1384
rect 5452 -1480 5772 -1448
rect 5452 -1486 5664 -1480
rect 4826 -1520 5374 -1492
rect 5140 -4080 5374 -1520
rect 5650 -1574 5664 -1486
rect 5654 -1594 5664 -1574
rect 5760 -1574 5772 -1480
rect 5760 -1594 5770 -1574
rect 5654 -1599 5770 -1594
rect 7050 -1666 7276 -1034
rect 7064 -1962 7276 -1666
rect 7050 -2356 7276 -1962
rect 7014 -2366 7522 -2356
rect 7014 -2368 7558 -2366
rect 7656 -2368 7766 -2364
rect 7014 -2478 7766 -2368
rect 7050 -2484 7766 -2478
rect 7050 -2488 7558 -2484
rect 7656 -2500 7766 -2484
rect 5138 -4086 5374 -4080
rect 5138 -4160 5372 -4086
rect 5132 -4192 5378 -4160
rect 5132 -4296 5148 -4192
rect 5364 -4296 5378 -4192
rect 5132 -4310 5378 -4296
<< via3 >>
rect 6790 -444 6954 -302
rect 8868 -464 9068 -312
rect 9554 -296 9686 -292
rect 9554 -406 9686 -296
rect 6478 -732 6640 -600
rect 9202 -752 9384 -582
rect 9688 -766 9760 -602
rect 9760 -766 9810 -602
rect 9688 -780 9810 -766
rect 6188 -1272 6320 -1172
rect 6188 -1282 6320 -1272
<< metal4 >>
rect 9734 -186 9735 -180
rect 6752 -282 6990 -258
rect 5548 -302 6998 -282
rect 5548 -444 6790 -302
rect 6954 -444 6998 -302
rect 5548 -450 6998 -444
rect 6440 -600 6678 -546
rect 6440 -732 6478 -600
rect 6640 -732 6678 -600
rect 6440 -792 6678 -732
rect 6752 -816 6990 -450
rect 7836 -812 8006 -218
rect 8850 -312 9086 -222
rect 9176 -232 9416 -190
rect 8850 -464 8868 -312
rect 9068 -464 9086 -312
rect 8850 -482 9086 -464
rect 9174 -582 9416 -232
rect 9484 -292 9734 -194
rect 9484 -406 9554 -292
rect 9686 -406 9734 -292
rect 9484 -422 9734 -406
rect 9486 -468 9734 -422
rect 9174 -752 9202 -582
rect 9384 -734 9416 -582
rect 9672 -602 9840 -576
rect 9384 -752 9414 -734
rect 9174 -776 9414 -752
rect 9672 -780 9688 -602
rect 9810 -780 9840 -602
rect 6187 -1172 6321 -1171
rect 6187 -1282 6188 -1172
rect 6320 -1282 6321 -1172
rect 9672 -1184 9840 -780
rect 6187 -1283 6321 -1282
rect 7944 -1358 9840 -1184
rect 9672 -1368 9840 -1358
use tt_asw_3v3  x1
timestamp 1731231864
transform 1 0 6104 0 1 -5137
box 0 0 3612 4352
use tt_asw_3v3  x2
timestamp 1731231864
transform -1 0 9755 0 -1 4116
box 0 0 3612 4352
use sky130_fd_sc_hd__inv_1  x3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731231864
transform -1 0 5218 0 1 -2556
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  x4 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1731231864
transform 0 1 5022 1 0 -1864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1731231864
transform 0 1 5002 1 0 -4138
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  x6
timestamp 1731231864
transform 0 1 5008 1 0 -3818
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1731231864
transform -1 0 5562 0 1 -2556
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x8
timestamp 1731231864
transform -1 0 5250 0 1 -3378
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1731231864
transform -1 0 5582 0 1 -3376
box -38 -48 314 592
<< labels >>
flabel metal1 5858 -454 6058 -254 0 FreeSans 256 0 0 0 VDDA
port 1 nsew
flabel metal1 9966 -772 10166 -572 0 FreeSans 256 0 0 0 VOUT
port 4 nsew
flabel metal1 5154 -1528 5354 -1328 0 FreeSans 256 0 0 0 Cin
port 2 nsew
flabel metal1 5540 -1308 5740 -1108 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 5536 -758 5736 -558 0 FreeSans 256 0 0 0 GND
port 0 nsew
<< end >>
