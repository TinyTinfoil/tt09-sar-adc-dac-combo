VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_veswaranandam_saradc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_veswaranandam_saradc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.330 77.750 97.330 77.830 ;
        RECT 75.440 71.370 97.330 77.750 ;
        RECT 71.420 71.330 101.250 71.370 ;
        RECT 71.420 67.390 101.330 71.330 ;
        RECT 71.440 67.330 101.330 67.390 ;
        RECT 71.440 67.250 100.370 67.330 ;
        RECT 75.440 66.830 100.370 67.250 ;
        RECT 75.440 66.750 86.440 66.830 ;
        RECT 96.330 61.690 100.370 66.830 ;
        RECT 96.300 57.650 100.400 61.690 ;
        RECT 89.950 21.545 94.650 21.550 ;
        RECT 89.775 16.855 94.825 21.545 ;
        RECT 89.950 8.030 94.650 16.855 ;
        RECT 89.950 3.330 136.750 8.030 ;
      LAYER met4 ;
        RECT 96.325 61.690 100.375 61.695 ;
        RECT 90.130 57.650 100.375 61.690 ;
        RECT 90.130 43.990 94.170 57.650 ;
        RECT 96.325 57.645 100.375 57.650 ;
        RECT 89.800 16.850 94.800 43.990 ;
        RECT 132.390 1.000 137.030 8.010 ;
        RECT 132.390 0.690 137.070 1.000 ;
        RECT 136.170 0.000 137.070 0.690 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 16.270 187.975 16.960 188.275 ;
        RECT 16.490 187.760 16.730 187.975 ;
        RECT 16.485 187.410 16.735 187.760 ;
        RECT 16.385 175.555 16.625 175.745 ;
        RECT 16.385 175.415 16.630 175.555 ;
        RECT 16.390 174.905 16.630 175.415 ;
        RECT 15.940 174.225 17.220 174.905 ;
      LAYER met1 ;
        RECT 16.070 188.145 17.070 189.145 ;
        RECT 16.310 188.005 16.900 188.145 ;
        RECT 15.990 174.255 17.180 174.885 ;
      LAYER met2 ;
        RECT 16.160 188.245 16.980 188.955 ;
        RECT 15.990 174.255 17.180 174.885 ;
      LAYER met3 ;
        RECT 14.320 217.560 15.210 217.570 ;
        RECT 122.380 217.560 123.200 224.130 ;
        RECT 14.320 216.520 123.310 217.560 ;
        RECT 14.320 189.195 15.210 216.520 ;
        RECT 14.320 189.175 17.160 189.195 ;
        RECT 14.320 188.185 17.170 189.175 ;
        RECT 14.320 188.150 15.210 188.185 ;
        RECT 16.000 175.385 17.170 188.185 ;
        RECT 15.990 175.355 17.170 175.385 ;
        RECT 15.990 174.985 17.160 175.355 ;
        RECT 15.960 174.235 17.190 174.985 ;
      LAYER met4 ;
        RECT 122.670 225.060 122.970 225.760 ;
        RECT 122.380 221.680 123.210 225.060 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 126.110 187.975 126.800 188.275 ;
        RECT 126.340 187.760 126.580 187.975 ;
        RECT 126.335 187.410 126.585 187.760 ;
        RECT 126.445 175.555 126.685 175.745 ;
        RECT 126.440 175.415 126.685 175.555 ;
        RECT 126.440 174.905 126.680 175.415 ;
        RECT 125.850 174.225 127.130 174.905 ;
      LAYER met1 ;
        RECT 126.000 188.145 127.000 189.145 ;
        RECT 126.170 188.005 126.760 188.145 ;
        RECT 125.890 174.255 127.080 174.885 ;
      LAYER met2 ;
        RECT 119.705 219.345 120.715 219.390 ;
        RECT 127.655 219.345 128.615 219.365 ;
        RECT 119.705 218.335 128.640 219.345 ;
        RECT 119.705 218.290 120.715 218.335 ;
        RECT 127.655 218.315 128.615 218.335 ;
        RECT 126.090 188.245 126.910 188.955 ;
        RECT 125.890 174.255 127.080 174.885 ;
      LAYER met3 ;
        RECT 119.630 221.745 120.440 224.210 ;
        RECT 119.630 221.640 120.715 221.745 ;
        RECT 119.620 220.050 120.715 221.640 ;
        RECT 119.490 219.370 120.715 220.050 ;
        RECT 119.490 218.310 120.740 219.370 ;
        RECT 119.490 218.120 120.130 218.310 ;
        RECT 127.630 189.195 128.640 219.415 ;
        RECT 125.910 189.175 128.640 189.195 ;
        RECT 125.900 188.185 128.640 189.175 ;
        RECT 125.900 175.385 127.070 188.185 ;
        RECT 125.900 175.355 127.080 175.385 ;
        RECT 125.910 174.985 127.080 175.355 ;
        RECT 125.880 174.235 127.110 174.985 ;
      LAYER met4 ;
        RECT 119.910 225.190 120.210 225.760 ;
        RECT 119.630 221.720 120.430 225.190 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 126.110 138.405 126.800 138.705 ;
        RECT 126.340 138.190 126.580 138.405 ;
        RECT 126.335 137.840 126.585 138.190 ;
        RECT 126.445 125.985 126.685 126.175 ;
        RECT 126.440 125.845 126.685 125.985 ;
        RECT 126.440 125.335 126.680 125.845 ;
        RECT 125.850 124.655 127.130 125.335 ;
      LAYER met1 ;
        RECT 126.000 138.575 127.000 139.575 ;
        RECT 126.170 138.435 126.760 138.575 ;
        RECT 125.890 124.685 127.080 125.315 ;
      LAYER met2 ;
        RECT 116.735 221.125 117.745 221.170 ;
        RECT 129.750 221.125 130.710 221.145 ;
        RECT 116.735 220.115 130.735 221.125 ;
        RECT 116.735 220.070 117.745 220.115 ;
        RECT 129.750 220.095 130.710 220.115 ;
        RECT 126.090 138.675 126.910 139.385 ;
        RECT 125.890 124.685 127.080 125.315 ;
      LAYER met3 ;
        RECT 116.800 223.340 117.650 224.360 ;
        RECT 116.760 222.150 117.800 223.340 ;
        RECT 116.760 222.065 117.900 222.150 ;
        RECT 116.735 221.150 117.900 222.065 ;
        RECT 116.710 221.140 117.900 221.150 ;
        RECT 116.710 220.090 117.770 221.140 ;
        RECT 129.725 220.115 133.705 221.125 ;
        RECT 132.695 170.645 133.705 220.115 ;
        RECT 127.630 169.635 133.705 170.645 ;
        RECT 127.630 139.625 128.640 169.635 ;
        RECT 125.910 139.605 128.640 139.625 ;
        RECT 125.900 138.615 128.640 139.605 ;
        RECT 125.900 125.815 127.070 138.615 ;
        RECT 125.900 125.785 127.080 125.815 ;
        RECT 125.910 125.415 127.080 125.785 ;
        RECT 125.880 124.665 127.110 125.415 ;
      LAYER met4 ;
        RECT 117.150 224.980 117.450 225.760 ;
        RECT 116.840 224.180 117.610 224.980 ;
        RECT 116.830 222.260 117.620 224.180 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 16.930 90.175 17.620 90.475 ;
        RECT 17.150 89.960 17.390 90.175 ;
        RECT 17.145 89.610 17.395 89.960 ;
        RECT 17.045 77.755 17.285 77.945 ;
        RECT 17.045 77.615 17.290 77.755 ;
        RECT 17.050 77.105 17.290 77.615 ;
        RECT 16.600 76.425 17.880 77.105 ;
      LAYER met1 ;
        RECT 16.730 90.345 17.730 91.345 ;
        RECT 16.970 90.205 17.560 90.345 ;
        RECT 16.650 76.455 17.840 77.085 ;
      LAYER met2 ;
        RECT 61.170 218.645 62.270 219.655 ;
        RECT 61.215 174.985 62.225 218.645 ;
        RECT 53.875 173.975 62.225 174.985 ;
        RECT 15.115 119.685 16.075 119.705 ;
        RECT 53.875 119.685 54.885 173.975 ;
        RECT 15.090 118.675 54.885 119.685 ;
        RECT 15.115 118.655 16.075 118.675 ;
        RECT 16.820 90.445 17.640 91.155 ;
        RECT 16.650 76.455 17.840 77.085 ;
      LAYER met3 ;
        RECT 113.990 223.445 114.840 224.420 ;
        RECT 113.855 223.310 114.865 223.445 ;
        RECT 113.855 221.320 114.930 223.310 ;
        RECT 61.190 219.655 62.250 219.680 ;
        RECT 113.855 219.655 114.865 221.320 ;
        RECT 61.190 218.645 114.865 219.655 ;
        RECT 61.190 218.620 62.250 218.645 ;
        RECT 15.090 91.395 16.100 119.685 ;
        RECT 15.090 91.375 17.820 91.395 ;
        RECT 15.090 90.385 17.830 91.375 ;
        RECT 16.660 77.585 17.830 90.385 ;
        RECT 16.650 77.555 17.830 77.585 ;
        RECT 16.650 77.185 17.820 77.555 ;
        RECT 16.620 76.435 17.850 77.185 ;
      LAYER met4 ;
        RECT 114.390 225.050 114.690 225.760 ;
        RECT 114.020 224.240 114.790 225.050 ;
        RECT 114.020 222.320 114.810 224.240 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 16.270 138.405 16.960 138.705 ;
        RECT 16.490 138.190 16.730 138.405 ;
        RECT 16.485 137.840 16.735 138.190 ;
        RECT 16.385 125.985 16.625 126.175 ;
        RECT 16.385 125.845 16.630 125.985 ;
        RECT 16.390 125.335 16.630 125.845 ;
        RECT 15.940 124.655 17.220 125.335 ;
      LAYER met1 ;
        RECT 16.070 138.575 17.070 139.575 ;
        RECT 16.310 138.435 16.900 138.575 ;
        RECT 15.990 124.685 17.180 125.315 ;
      LAYER met2 ;
        RECT 56.895 220.680 58.160 221.855 ;
        RECT 56.940 180.255 58.115 220.680 ;
        RECT 39.735 179.080 58.115 180.255 ;
        RECT 39.735 168.455 40.910 179.080 ;
        RECT 39.720 167.345 40.920 168.455 ;
        RECT 39.735 167.315 40.910 167.345 ;
        RECT 16.160 138.675 16.980 139.385 ;
        RECT 15.990 124.685 17.180 125.315 ;
      LAYER met3 ;
        RECT 111.390 223.230 112.240 224.430 ;
        RECT 111.260 222.725 112.300 223.230 ;
        RECT 56.915 221.855 58.140 221.880 ;
        RECT 111.260 221.855 112.495 222.725 ;
        RECT 56.915 220.680 112.495 221.855 ;
        RECT 56.915 220.655 58.140 220.680 ;
        RECT 11.480 167.320 41.590 168.480 ;
        RECT 11.480 139.625 12.640 167.320 ;
        RECT 11.480 139.605 17.160 139.625 ;
        RECT 11.480 138.615 17.170 139.605 ;
        RECT 11.480 138.540 12.640 138.615 ;
        RECT 16.000 125.815 17.170 138.615 ;
        RECT 15.990 125.785 17.170 125.815 ;
        RECT 15.990 125.415 17.160 125.785 ;
        RECT 15.960 124.665 17.190 125.415 ;
      LAYER met4 ;
        RECT 111.630 225.050 111.930 225.760 ;
        RECT 111.410 224.040 112.210 225.050 ;
        RECT 111.420 222.330 112.210 224.040 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 126.110 89.505 126.800 89.805 ;
        RECT 126.340 89.290 126.580 89.505 ;
        RECT 126.335 88.940 126.585 89.290 ;
        RECT 126.445 77.085 126.685 77.275 ;
        RECT 126.440 76.945 126.685 77.085 ;
        RECT 126.440 76.435 126.680 76.945 ;
        RECT 125.850 75.755 127.130 76.435 ;
      LAYER met1 ;
        RECT 126.000 89.675 127.000 90.675 ;
        RECT 126.170 89.535 126.760 89.675 ;
        RECT 125.890 75.785 127.080 76.415 ;
      LAYER met2 ;
        RECT 108.395 218.795 109.405 224.100 ;
        RECT 100.535 217.785 109.405 218.795 ;
        RECT 100.535 204.955 101.545 217.785 ;
        RECT 83.105 203.945 101.545 204.955 ;
        RECT 83.105 119.385 84.115 203.945 ;
        RECT 123.760 119.385 124.720 119.405 ;
        RECT 83.105 118.375 124.745 119.385 ;
        RECT 123.760 118.355 124.720 118.375 ;
        RECT 126.090 89.775 126.910 90.485 ;
        RECT 125.890 75.785 127.080 76.415 ;
      LAYER met3 ;
        RECT 108.395 224.080 109.405 224.685 ;
        RECT 108.370 223.020 109.430 224.080 ;
        RECT 123.735 118.375 128.640 119.385 ;
        RECT 127.630 90.725 128.640 118.375 ;
        RECT 125.910 90.705 128.640 90.725 ;
        RECT 125.900 89.715 128.640 90.705 ;
        RECT 125.900 76.915 127.070 89.715 ;
        RECT 125.900 76.885 127.080 76.915 ;
        RECT 125.910 76.515 127.080 76.885 ;
        RECT 125.880 75.765 127.110 76.515 ;
      LAYER met4 ;
        RECT 108.395 224.660 109.405 225.845 ;
        RECT 108.390 223.640 109.410 224.660 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 125.450 39.605 126.140 39.905 ;
        RECT 125.680 39.390 125.920 39.605 ;
        RECT 125.675 39.040 125.925 39.390 ;
        RECT 125.785 27.185 126.025 27.375 ;
        RECT 125.780 27.045 126.025 27.185 ;
        RECT 125.780 26.535 126.020 27.045 ;
        RECT 125.190 25.855 126.470 26.535 ;
      LAYER met1 ;
        RECT 125.340 39.775 126.340 40.775 ;
        RECT 125.510 39.635 126.100 39.775 ;
        RECT 125.230 25.885 126.420 26.515 ;
      LAYER met2 ;
        RECT 75.450 222.875 76.550 223.885 ;
        RECT 75.495 109.515 76.505 222.875 ;
        RECT 75.495 108.505 83.565 109.515 ;
        RECT 82.555 70.235 83.565 108.505 ;
        RECT 126.995 70.235 127.955 70.255 ;
        RECT 82.555 69.225 127.980 70.235 ;
        RECT 126.995 69.205 127.955 69.225 ;
        RECT 125.430 39.875 126.250 40.585 ;
        RECT 125.230 25.885 126.420 26.515 ;
      LAYER met3 ;
        RECT 75.470 223.885 76.530 223.910 ;
        RECT 75.470 222.875 79.315 223.885 ;
        RECT 75.470 222.850 76.530 222.875 ;
        RECT 126.970 40.825 127.980 70.235 ;
        RECT 125.250 40.805 127.980 40.825 ;
        RECT 125.240 39.815 127.980 40.805 ;
        RECT 125.240 27.015 126.410 39.815 ;
        RECT 125.240 26.985 126.420 27.015 ;
        RECT 125.250 26.615 126.420 26.985 ;
        RECT 125.220 25.865 126.450 26.615 ;
      LAYER met4 ;
        RECT 106.110 225.545 106.410 225.760 ;
        RECT 78.270 223.885 79.290 223.890 ;
        RECT 78.270 222.875 100.085 223.885 ;
        RECT 78.270 222.870 79.290 222.875 ;
        RECT 99.075 220.485 100.085 222.875 ;
        RECT 105.525 220.485 106.535 225.545 ;
        RECT 99.075 219.475 106.535 220.485 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 16.600 39.605 17.290 39.905 ;
        RECT 16.820 39.390 17.060 39.605 ;
        RECT 16.815 39.040 17.065 39.390 ;
        RECT 16.715 27.185 16.955 27.375 ;
        RECT 16.715 27.045 16.960 27.185 ;
        RECT 16.720 26.535 16.960 27.045 ;
        RECT 16.270 25.855 17.550 26.535 ;
      LAYER met1 ;
        RECT 102.715 219.465 103.725 223.845 ;
        RECT 54.565 218.455 103.725 219.465 ;
        RECT 20.615 70.345 21.625 70.375 ;
        RECT 54.565 70.345 55.575 218.455 ;
        RECT 20.615 69.335 55.575 70.345 ;
        RECT 20.615 69.305 21.625 69.335 ;
        RECT 16.400 39.775 17.400 40.775 ;
        RECT 16.640 39.635 17.230 39.775 ;
        RECT 16.320 25.885 17.510 26.515 ;
      LAYER met2 ;
        RECT 102.715 223.815 103.725 224.500 ;
        RECT 102.685 222.805 103.755 223.815 ;
        RECT 14.760 70.320 21.655 70.345 ;
        RECT 14.740 69.360 21.655 70.320 ;
        RECT 14.760 69.335 21.655 69.360 ;
        RECT 16.490 39.875 17.310 40.585 ;
        RECT 16.320 25.885 17.510 26.515 ;
      LAYER met3 ;
        RECT 102.715 224.480 103.725 225.075 ;
        RECT 102.690 223.420 103.750 224.480 ;
        RECT 14.760 40.825 15.770 70.345 ;
        RECT 14.760 40.805 17.490 40.825 ;
        RECT 14.760 39.815 17.500 40.805 ;
        RECT 16.330 27.015 17.500 39.815 ;
        RECT 16.320 26.985 17.500 27.015 ;
        RECT 16.320 26.615 17.490 26.985 ;
        RECT 16.290 25.865 17.520 26.615 ;
      LAYER met4 ;
        RECT 102.715 225.050 103.725 225.785 ;
        RECT 102.710 224.030 103.730 225.050 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 37.525 195.005 38.885 196.365 ;
        RECT 104.185 195.005 105.545 196.365 ;
        RECT 21.010 190.100 22.370 191.460 ;
        RECT 120.700 190.100 122.060 191.460 ;
        RECT 37.525 145.435 38.885 146.795 ;
        RECT 104.185 145.435 105.545 146.795 ;
        RECT 21.010 140.530 22.370 141.890 ;
        RECT 120.700 140.530 122.060 141.890 ;
        RECT 38.185 97.205 39.545 98.565 ;
        RECT 104.185 96.535 105.545 97.895 ;
        RECT 21.670 92.300 23.030 93.660 ;
        RECT 120.700 91.630 122.060 92.990 ;
        RECT 37.855 46.635 39.215 47.995 ;
        RECT 103.525 46.635 104.885 47.995 ;
        RECT 21.340 41.730 22.700 43.090 ;
        RECT 120.040 41.730 121.400 43.090 ;
      LAYER li1 ;
        RECT 37.745 195.115 38.665 195.785 ;
        RECT 104.405 195.115 105.325 195.785 ;
        RECT 21.230 190.680 22.150 191.350 ;
        RECT 120.920 190.680 121.840 191.350 ;
        RECT 18.045 187.750 18.215 187.845 ;
        RECT 16.905 187.420 18.215 187.750 ;
        RECT 18.045 186.465 18.215 187.420 ;
        RECT 124.855 187.750 125.025 187.845 ;
        RECT 124.855 187.420 126.165 187.750 ;
        RECT 124.855 186.465 125.025 187.420 ;
        RECT 15.010 185.640 16.390 185.810 ;
        RECT 16.730 185.640 18.110 185.810 ;
        RECT 124.960 185.640 126.340 185.810 ;
        RECT 126.680 185.640 128.060 185.810 ;
        RECT 15.840 184.500 16.050 185.640 ;
        RECT 17.560 184.500 17.770 185.640 ;
        RECT 125.300 184.500 125.510 185.640 ;
        RECT 127.020 184.500 127.230 185.640 ;
        RECT 15.170 181.530 16.550 181.700 ;
        RECT 16.830 181.540 18.210 181.710 ;
        RECT 124.860 181.540 126.240 181.710 ;
        RECT 16.000 180.390 16.210 181.530 ;
        RECT 17.660 180.400 17.870 181.540 ;
        RECT 125.200 180.400 125.410 181.540 ;
        RECT 126.520 181.530 127.900 181.700 ;
        RECT 126.860 180.390 127.070 181.530 ;
        RECT 17.975 177.980 18.145 178.075 ;
        RECT 16.835 177.650 18.145 177.980 ;
        RECT 17.975 176.695 18.145 177.650 ;
        RECT 124.925 177.980 125.095 178.075 ;
        RECT 124.925 177.650 126.235 177.980 ;
        RECT 124.925 176.695 125.095 177.650 ;
        RECT 17.945 175.645 18.115 176.475 ;
        RECT 16.805 175.435 18.115 175.645 ;
        RECT 17.945 175.095 18.115 175.435 ;
        RECT 124.955 175.645 125.125 176.475 ;
        RECT 124.955 175.435 126.265 175.645 ;
        RECT 124.955 175.095 125.125 175.435 ;
        RECT 37.745 145.545 38.665 146.215 ;
        RECT 104.405 145.545 105.325 146.215 ;
        RECT 21.230 141.110 22.150 141.780 ;
        RECT 120.920 141.110 121.840 141.780 ;
        RECT 18.045 138.180 18.215 138.275 ;
        RECT 16.905 137.850 18.215 138.180 ;
        RECT 18.045 136.895 18.215 137.850 ;
        RECT 124.855 138.180 125.025 138.275 ;
        RECT 124.855 137.850 126.165 138.180 ;
        RECT 124.855 136.895 125.025 137.850 ;
        RECT 15.010 136.070 16.390 136.240 ;
        RECT 16.730 136.070 18.110 136.240 ;
        RECT 124.960 136.070 126.340 136.240 ;
        RECT 126.680 136.070 128.060 136.240 ;
        RECT 15.840 134.930 16.050 136.070 ;
        RECT 17.560 134.930 17.770 136.070 ;
        RECT 125.300 134.930 125.510 136.070 ;
        RECT 127.020 134.930 127.230 136.070 ;
        RECT 15.170 131.960 16.550 132.130 ;
        RECT 16.830 131.970 18.210 132.140 ;
        RECT 124.860 131.970 126.240 132.140 ;
        RECT 16.000 130.820 16.210 131.960 ;
        RECT 17.660 130.830 17.870 131.970 ;
        RECT 125.200 130.830 125.410 131.970 ;
        RECT 126.520 131.960 127.900 132.130 ;
        RECT 126.860 130.820 127.070 131.960 ;
        RECT 17.975 128.410 18.145 128.505 ;
        RECT 16.835 128.080 18.145 128.410 ;
        RECT 17.975 127.125 18.145 128.080 ;
        RECT 124.925 128.410 125.095 128.505 ;
        RECT 124.925 128.080 126.235 128.410 ;
        RECT 124.925 127.125 125.095 128.080 ;
        RECT 17.945 126.075 18.115 126.905 ;
        RECT 16.805 125.865 18.115 126.075 ;
        RECT 17.945 125.525 18.115 125.865 ;
        RECT 124.955 126.075 125.125 126.905 ;
        RECT 124.955 125.865 126.265 126.075 ;
        RECT 124.955 125.525 125.125 125.865 ;
        RECT 38.405 97.315 39.325 97.985 ;
        RECT 104.405 96.645 105.325 97.315 ;
        RECT 21.890 92.880 22.810 93.550 ;
        RECT 120.920 92.210 121.840 92.880 ;
        RECT 18.705 89.950 18.875 90.045 ;
        RECT 17.565 89.620 18.875 89.950 ;
        RECT 18.705 88.665 18.875 89.620 ;
        RECT 124.855 89.280 125.025 89.375 ;
        RECT 124.855 88.950 126.165 89.280 ;
        RECT 15.670 87.840 17.050 88.010 ;
        RECT 17.390 87.840 18.770 88.010 ;
        RECT 124.855 87.995 125.025 88.950 ;
        RECT 16.500 86.700 16.710 87.840 ;
        RECT 18.220 86.700 18.430 87.840 ;
        RECT 124.960 87.170 126.340 87.340 ;
        RECT 126.680 87.170 128.060 87.340 ;
        RECT 125.300 86.030 125.510 87.170 ;
        RECT 127.020 86.030 127.230 87.170 ;
        RECT 15.830 83.730 17.210 83.900 ;
        RECT 17.490 83.740 18.870 83.910 ;
        RECT 16.660 82.590 16.870 83.730 ;
        RECT 18.320 82.600 18.530 83.740 ;
        RECT 124.860 83.070 126.240 83.240 ;
        RECT 125.200 81.930 125.410 83.070 ;
        RECT 126.520 83.060 127.900 83.230 ;
        RECT 126.860 81.920 127.070 83.060 ;
        RECT 18.635 80.180 18.805 80.275 ;
        RECT 17.495 79.850 18.805 80.180 ;
        RECT 18.635 78.895 18.805 79.850 ;
        RECT 124.925 79.510 125.095 79.605 ;
        RECT 124.925 79.180 126.235 79.510 ;
        RECT 18.605 77.845 18.775 78.675 ;
        RECT 124.925 78.225 125.095 79.180 ;
        RECT 17.465 77.635 18.775 77.845 ;
        RECT 18.605 77.295 18.775 77.635 ;
        RECT 124.955 77.175 125.125 78.005 ;
        RECT 124.955 76.965 126.265 77.175 ;
        RECT 124.955 76.625 125.125 76.965 ;
        RECT 38.075 46.745 38.995 47.415 ;
        RECT 103.745 46.745 104.665 47.415 ;
        RECT 21.560 42.310 22.480 42.980 ;
        RECT 120.260 42.310 121.180 42.980 ;
        RECT 18.375 39.380 18.545 39.475 ;
        RECT 17.235 39.050 18.545 39.380 ;
        RECT 18.375 38.095 18.545 39.050 ;
        RECT 124.195 39.380 124.365 39.475 ;
        RECT 124.195 39.050 125.505 39.380 ;
        RECT 124.195 38.095 124.365 39.050 ;
        RECT 15.340 37.270 16.720 37.440 ;
        RECT 17.060 37.270 18.440 37.440 ;
        RECT 124.300 37.270 125.680 37.440 ;
        RECT 126.020 37.270 127.400 37.440 ;
        RECT 16.170 36.130 16.380 37.270 ;
        RECT 17.890 36.130 18.100 37.270 ;
        RECT 124.640 36.130 124.850 37.270 ;
        RECT 126.360 36.130 126.570 37.270 ;
        RECT 15.500 33.160 16.880 33.330 ;
        RECT 17.160 33.170 18.540 33.340 ;
        RECT 124.200 33.170 125.580 33.340 ;
        RECT 16.330 32.020 16.540 33.160 ;
        RECT 17.990 32.030 18.200 33.170 ;
        RECT 124.540 32.030 124.750 33.170 ;
        RECT 125.860 33.160 127.240 33.330 ;
        RECT 126.200 32.020 126.410 33.160 ;
        RECT 18.305 29.610 18.475 29.705 ;
        RECT 17.165 29.280 18.475 29.610 ;
        RECT 18.305 28.325 18.475 29.280 ;
        RECT 124.265 29.610 124.435 29.705 ;
        RECT 124.265 29.280 125.575 29.610 ;
        RECT 124.265 28.325 124.435 29.280 ;
        RECT 18.275 27.275 18.445 28.105 ;
        RECT 17.135 27.065 18.445 27.275 ;
        RECT 18.275 26.725 18.445 27.065 ;
        RECT 124.295 27.275 124.465 28.105 ;
        RECT 124.295 27.065 125.605 27.275 ;
        RECT 124.295 26.725 124.465 27.065 ;
      LAYER met1 ;
        RECT 37.745 195.115 38.665 195.715 ;
        RECT 104.405 195.115 105.325 195.715 ;
        RECT 21.230 190.750 22.150 191.350 ;
        RECT 120.920 190.750 121.840 191.350 ;
        RECT 17.870 190.245 18.380 190.255 ;
        RECT 124.690 190.245 125.200 190.255 ;
        RECT 17.870 189.245 19.000 190.245 ;
        RECT 124.070 189.245 125.200 190.245 ;
        RECT 17.870 189.125 18.410 189.245 ;
        RECT 17.900 188.315 18.410 189.125 ;
        RECT 124.660 189.125 125.200 189.245 ;
        RECT 124.660 188.315 125.170 189.125 ;
        RECT 17.900 187.845 18.390 188.315 ;
        RECT 17.890 187.825 18.390 187.845 ;
        RECT 124.680 187.845 125.170 188.315 ;
        RECT 124.680 187.825 125.180 187.845 ;
        RECT 17.890 186.465 18.370 187.825 ;
        RECT 124.700 186.465 125.180 187.825 ;
        RECT 17.890 185.965 18.360 186.465 ;
        RECT 15.010 185.935 18.360 185.965 ;
        RECT 124.710 185.965 125.180 186.465 ;
        RECT 124.710 185.935 128.060 185.965 ;
        RECT 15.010 185.485 19.050 185.935 ;
        RECT 17.890 185.475 19.050 185.485 ;
        RECT 18.270 185.465 19.050 185.475 ;
        RECT 124.020 185.485 128.060 185.935 ;
        RECT 124.020 185.475 125.180 185.485 ;
        RECT 124.020 185.465 124.800 185.475 ;
        RECT 18.350 182.005 19.040 185.465 ;
        RECT 124.030 182.005 124.720 185.465 ;
        RECT 18.350 181.865 19.190 182.005 ;
        RECT 123.880 181.865 124.720 182.005 ;
        RECT 16.450 181.855 18.210 181.865 ;
        RECT 18.350 181.855 21.320 181.865 ;
        RECT 121.750 181.855 124.720 181.865 ;
        RECT 124.860 181.855 126.620 181.865 ;
        RECT 15.170 181.395 21.770 181.855 ;
        RECT 15.170 181.385 18.210 181.395 ;
        RECT 15.170 181.375 16.870 181.385 ;
        RECT 21.230 180.585 21.770 181.395 ;
        RECT 21.210 180.465 21.770 180.585 ;
        RECT 121.300 181.395 127.900 181.855 ;
        RECT 121.300 180.585 121.840 181.395 ;
        RECT 124.860 181.385 127.900 181.395 ;
        RECT 126.200 181.375 127.900 181.385 ;
        RECT 121.300 180.465 121.860 180.585 ;
        RECT 21.210 178.105 21.750 180.465 ;
        RECT 19.900 178.085 21.750 178.105 ;
        RECT 19.360 178.075 21.750 178.085 ;
        RECT 17.820 178.055 21.750 178.075 ;
        RECT 121.320 178.105 121.860 180.465 ;
        RECT 121.320 178.085 123.170 178.105 ;
        RECT 121.320 178.075 123.710 178.085 ;
        RECT 121.320 178.055 125.250 178.075 ;
        RECT 17.820 177.635 21.760 178.055 ;
        RECT 17.820 176.745 18.300 177.635 ;
        RECT 18.940 177.615 21.760 177.635 ;
        RECT 121.310 177.635 125.250 178.055 ;
        RECT 121.310 177.615 124.130 177.635 ;
        RECT 19.360 177.605 21.080 177.615 ;
        RECT 121.990 177.605 123.710 177.615 ;
        RECT 17.810 176.695 18.300 176.745 ;
        RECT 124.770 176.745 125.250 177.635 ;
        RECT 124.770 176.695 125.260 176.745 ;
        RECT 17.810 176.475 18.290 176.695 ;
        RECT 17.790 176.415 18.290 176.475 ;
        RECT 124.780 176.475 125.260 176.695 ;
        RECT 124.780 176.415 125.280 176.475 ;
        RECT 17.790 175.095 18.270 176.415 ;
        RECT 124.800 175.095 125.280 176.415 ;
        RECT 37.745 145.545 38.665 146.145 ;
        RECT 104.405 145.545 105.325 146.145 ;
        RECT 21.230 141.180 22.150 141.780 ;
        RECT 120.920 141.180 121.840 141.780 ;
        RECT 17.870 140.675 18.380 140.685 ;
        RECT 124.690 140.675 125.200 140.685 ;
        RECT 17.870 139.675 19.000 140.675 ;
        RECT 124.070 139.675 125.200 140.675 ;
        RECT 17.870 139.555 18.410 139.675 ;
        RECT 17.900 138.745 18.410 139.555 ;
        RECT 124.660 139.555 125.200 139.675 ;
        RECT 124.660 138.745 125.170 139.555 ;
        RECT 17.900 138.275 18.390 138.745 ;
        RECT 17.890 138.255 18.390 138.275 ;
        RECT 124.680 138.275 125.170 138.745 ;
        RECT 124.680 138.255 125.180 138.275 ;
        RECT 17.890 136.895 18.370 138.255 ;
        RECT 124.700 136.895 125.180 138.255 ;
        RECT 17.890 136.395 18.360 136.895 ;
        RECT 15.010 136.365 18.360 136.395 ;
        RECT 124.710 136.395 125.180 136.895 ;
        RECT 124.710 136.365 128.060 136.395 ;
        RECT 15.010 135.915 19.050 136.365 ;
        RECT 17.890 135.905 19.050 135.915 ;
        RECT 18.270 135.895 19.050 135.905 ;
        RECT 124.020 135.915 128.060 136.365 ;
        RECT 124.020 135.905 125.180 135.915 ;
        RECT 124.020 135.895 124.800 135.905 ;
        RECT 18.350 132.435 19.040 135.895 ;
        RECT 124.030 132.435 124.720 135.895 ;
        RECT 18.350 132.295 19.190 132.435 ;
        RECT 123.880 132.295 124.720 132.435 ;
        RECT 16.450 132.285 18.210 132.295 ;
        RECT 18.350 132.285 21.320 132.295 ;
        RECT 121.750 132.285 124.720 132.295 ;
        RECT 124.860 132.285 126.620 132.295 ;
        RECT 15.170 131.825 21.770 132.285 ;
        RECT 15.170 131.815 18.210 131.825 ;
        RECT 15.170 131.805 16.870 131.815 ;
        RECT 21.230 131.015 21.770 131.825 ;
        RECT 21.210 130.895 21.770 131.015 ;
        RECT 121.300 131.825 127.900 132.285 ;
        RECT 121.300 131.015 121.840 131.825 ;
        RECT 124.860 131.815 127.900 131.825 ;
        RECT 126.200 131.805 127.900 131.815 ;
        RECT 121.300 130.895 121.860 131.015 ;
        RECT 21.210 128.535 21.750 130.895 ;
        RECT 19.900 128.515 21.750 128.535 ;
        RECT 19.360 128.505 21.750 128.515 ;
        RECT 17.820 128.485 21.750 128.505 ;
        RECT 121.320 128.535 121.860 130.895 ;
        RECT 121.320 128.515 123.170 128.535 ;
        RECT 121.320 128.505 123.710 128.515 ;
        RECT 121.320 128.485 125.250 128.505 ;
        RECT 17.820 128.065 21.760 128.485 ;
        RECT 17.820 127.175 18.300 128.065 ;
        RECT 18.940 128.045 21.760 128.065 ;
        RECT 121.310 128.065 125.250 128.485 ;
        RECT 121.310 128.045 124.130 128.065 ;
        RECT 19.360 128.035 21.080 128.045 ;
        RECT 121.990 128.035 123.710 128.045 ;
        RECT 17.810 127.125 18.300 127.175 ;
        RECT 124.770 127.175 125.250 128.065 ;
        RECT 124.770 127.125 125.260 127.175 ;
        RECT 17.810 126.905 18.290 127.125 ;
        RECT 17.790 126.845 18.290 126.905 ;
        RECT 124.780 126.905 125.260 127.125 ;
        RECT 124.780 126.845 125.280 126.905 ;
        RECT 17.790 125.525 18.270 126.845 ;
        RECT 124.800 125.525 125.280 126.845 ;
        RECT 38.405 97.315 39.325 97.915 ;
        RECT 104.405 96.645 105.325 97.245 ;
        RECT 21.890 92.950 22.810 93.550 ;
        RECT 18.530 92.445 19.040 92.455 ;
        RECT 18.530 91.445 19.660 92.445 ;
        RECT 120.920 92.280 121.840 92.880 ;
        RECT 124.690 91.775 125.200 91.785 ;
        RECT 18.530 91.325 19.070 91.445 ;
        RECT 18.560 90.515 19.070 91.325 ;
        RECT 124.070 90.775 125.200 91.775 ;
        RECT 124.660 90.655 125.200 90.775 ;
        RECT 18.560 90.045 19.050 90.515 ;
        RECT 18.550 90.025 19.050 90.045 ;
        RECT 18.550 88.665 19.030 90.025 ;
        RECT 124.660 89.845 125.170 90.655 ;
        RECT 124.680 89.375 125.170 89.845 ;
        RECT 124.680 89.355 125.180 89.375 ;
        RECT 18.550 88.165 19.020 88.665 ;
        RECT 15.670 88.135 19.020 88.165 ;
        RECT 15.670 87.685 19.710 88.135 ;
        RECT 124.700 87.995 125.180 89.355 ;
        RECT 18.550 87.675 19.710 87.685 ;
        RECT 18.930 87.665 19.710 87.675 ;
        RECT 19.010 84.205 19.700 87.665 ;
        RECT 124.710 87.495 125.180 87.995 ;
        RECT 124.710 87.465 128.060 87.495 ;
        RECT 124.020 87.015 128.060 87.465 ;
        RECT 124.020 87.005 125.180 87.015 ;
        RECT 124.020 86.995 124.800 87.005 ;
        RECT 19.010 84.065 19.850 84.205 ;
        RECT 17.110 84.055 18.870 84.065 ;
        RECT 19.010 84.055 21.980 84.065 ;
        RECT 15.830 83.595 22.430 84.055 ;
        RECT 15.830 83.585 18.870 83.595 ;
        RECT 15.830 83.575 17.530 83.585 ;
        RECT 21.890 82.785 22.430 83.595 ;
        RECT 124.030 83.535 124.720 86.995 ;
        RECT 123.880 83.395 124.720 83.535 ;
        RECT 121.750 83.385 124.720 83.395 ;
        RECT 124.860 83.385 126.620 83.395 ;
        RECT 21.870 82.665 22.430 82.785 ;
        RECT 121.300 82.925 127.900 83.385 ;
        RECT 21.870 80.305 22.410 82.665 ;
        RECT 121.300 82.115 121.840 82.925 ;
        RECT 124.860 82.915 127.900 82.925 ;
        RECT 126.200 82.905 127.900 82.915 ;
        RECT 121.300 81.995 121.860 82.115 ;
        RECT 20.560 80.285 22.410 80.305 ;
        RECT 20.020 80.275 22.410 80.285 ;
        RECT 18.480 80.255 22.410 80.275 ;
        RECT 18.480 79.835 22.420 80.255 ;
        RECT 18.480 78.945 18.960 79.835 ;
        RECT 19.600 79.815 22.420 79.835 ;
        RECT 20.020 79.805 21.740 79.815 ;
        RECT 121.320 79.635 121.860 81.995 ;
        RECT 121.320 79.615 123.170 79.635 ;
        RECT 121.320 79.605 123.710 79.615 ;
        RECT 121.320 79.585 125.250 79.605 ;
        RECT 121.310 79.165 125.250 79.585 ;
        RECT 121.310 79.145 124.130 79.165 ;
        RECT 121.990 79.135 123.710 79.145 ;
        RECT 18.470 78.895 18.960 78.945 ;
        RECT 18.470 78.675 18.950 78.895 ;
        RECT 18.450 78.615 18.950 78.675 ;
        RECT 18.450 77.295 18.930 78.615 ;
        RECT 124.770 78.275 125.250 79.165 ;
        RECT 124.770 78.225 125.260 78.275 ;
        RECT 124.780 78.005 125.260 78.225 ;
        RECT 124.780 77.945 125.280 78.005 ;
        RECT 124.800 76.625 125.280 77.945 ;
        RECT 38.075 46.745 38.995 47.345 ;
        RECT 103.745 46.745 104.665 47.345 ;
        RECT 21.560 42.380 22.480 42.980 ;
        RECT 120.260 42.380 121.180 42.980 ;
        RECT 18.200 41.875 18.710 41.885 ;
        RECT 124.030 41.875 124.540 41.885 ;
        RECT 18.200 40.875 19.330 41.875 ;
        RECT 123.410 40.875 124.540 41.875 ;
        RECT 18.200 40.755 18.740 40.875 ;
        RECT 18.230 39.945 18.740 40.755 ;
        RECT 124.000 40.755 124.540 40.875 ;
        RECT 124.000 39.945 124.510 40.755 ;
        RECT 18.230 39.475 18.720 39.945 ;
        RECT 18.220 39.455 18.720 39.475 ;
        RECT 124.020 39.475 124.510 39.945 ;
        RECT 124.020 39.455 124.520 39.475 ;
        RECT 18.220 38.095 18.700 39.455 ;
        RECT 124.040 38.095 124.520 39.455 ;
        RECT 18.220 37.595 18.690 38.095 ;
        RECT 15.340 37.565 18.690 37.595 ;
        RECT 124.050 37.595 124.520 38.095 ;
        RECT 124.050 37.565 127.400 37.595 ;
        RECT 15.340 37.115 19.380 37.565 ;
        RECT 18.220 37.105 19.380 37.115 ;
        RECT 18.600 37.095 19.380 37.105 ;
        RECT 123.360 37.115 127.400 37.565 ;
        RECT 123.360 37.105 124.520 37.115 ;
        RECT 123.360 37.095 124.140 37.105 ;
        RECT 18.680 33.635 19.370 37.095 ;
        RECT 123.370 33.635 124.060 37.095 ;
        RECT 18.680 33.495 19.520 33.635 ;
        RECT 123.220 33.495 124.060 33.635 ;
        RECT 16.780 33.485 18.540 33.495 ;
        RECT 18.680 33.485 21.650 33.495 ;
        RECT 121.090 33.485 124.060 33.495 ;
        RECT 124.200 33.485 125.960 33.495 ;
        RECT 15.500 33.025 22.100 33.485 ;
        RECT 15.500 33.015 18.540 33.025 ;
        RECT 15.500 33.005 17.200 33.015 ;
        RECT 21.560 32.215 22.100 33.025 ;
        RECT 21.540 32.095 22.100 32.215 ;
        RECT 120.640 33.025 127.240 33.485 ;
        RECT 120.640 32.215 121.180 33.025 ;
        RECT 124.200 33.015 127.240 33.025 ;
        RECT 125.540 33.005 127.240 33.015 ;
        RECT 120.640 32.095 121.200 32.215 ;
        RECT 21.540 29.735 22.080 32.095 ;
        RECT 20.230 29.715 22.080 29.735 ;
        RECT 19.690 29.705 22.080 29.715 ;
        RECT 18.150 29.685 22.080 29.705 ;
        RECT 120.660 29.735 121.200 32.095 ;
        RECT 120.660 29.715 122.510 29.735 ;
        RECT 120.660 29.705 123.050 29.715 ;
        RECT 120.660 29.685 124.590 29.705 ;
        RECT 18.150 29.265 22.090 29.685 ;
        RECT 18.150 28.375 18.630 29.265 ;
        RECT 19.270 29.245 22.090 29.265 ;
        RECT 120.650 29.265 124.590 29.685 ;
        RECT 120.650 29.245 123.470 29.265 ;
        RECT 19.690 29.235 21.410 29.245 ;
        RECT 121.330 29.235 123.050 29.245 ;
        RECT 18.140 28.325 18.630 28.375 ;
        RECT 124.110 28.375 124.590 29.265 ;
        RECT 124.110 28.325 124.600 28.375 ;
        RECT 18.140 28.105 18.620 28.325 ;
        RECT 18.120 28.045 18.620 28.105 ;
        RECT 124.120 28.105 124.600 28.325 ;
        RECT 124.120 28.045 124.620 28.105 ;
        RECT 18.120 26.725 18.600 28.045 ;
        RECT 124.140 26.725 124.620 28.045 ;
      LAYER met2 ;
        RECT 37.745 195.215 38.665 195.545 ;
        RECT 104.405 195.215 105.325 195.545 ;
        RECT 37.730 194.165 38.970 194.585 ;
        RECT 25.920 193.445 38.970 194.165 ;
        RECT 104.100 194.165 105.340 194.585 ;
        RECT 104.100 193.445 117.150 194.165 ;
        RECT 25.920 193.395 38.230 193.445 ;
        RECT 104.840 193.395 117.150 193.445 ;
        RECT 25.920 192.015 26.580 193.395 ;
        RECT 116.490 192.015 117.150 193.395 ;
        RECT 25.910 191.855 26.650 192.015 ;
        RECT 21.230 190.920 22.150 191.250 ;
        RECT 25.920 190.675 26.650 191.855 ;
        RECT 1.100 190.260 2.840 190.560 ;
        RECT 1.100 190.220 6.160 190.260 ;
        RECT 1.100 190.185 17.120 190.220 ;
        RECT 1.100 190.145 18.160 190.185 ;
        RECT 1.100 190.105 18.650 190.145 ;
        RECT 19.300 190.105 21.160 190.125 ;
        RECT 25.910 190.115 26.650 190.675 ;
        RECT 1.100 190.095 21.880 190.105 ;
        RECT 23.900 190.095 26.650 190.115 ;
        RECT 1.100 189.455 26.650 190.095 ;
        RECT 1.100 189.355 22.650 189.455 ;
        RECT 23.580 189.355 26.650 189.455 ;
        RECT 1.100 189.325 21.880 189.355 ;
        RECT 25.910 189.345 26.650 189.355 ;
        RECT 116.420 191.855 117.160 192.015 ;
        RECT 116.420 190.675 117.150 191.855 ;
        RECT 120.920 190.920 121.840 191.250 ;
        RECT 116.420 190.115 117.160 190.675 ;
        RECT 132.315 190.185 134.805 223.135 ;
        RECT 124.910 190.145 134.805 190.185 ;
        RECT 116.420 190.095 119.170 190.115 ;
        RECT 121.910 190.105 123.770 190.125 ;
        RECT 124.420 190.105 134.805 190.145 ;
        RECT 121.190 190.095 134.805 190.105 ;
        RECT 116.420 189.455 134.805 190.095 ;
        RECT 116.420 189.355 119.490 189.455 ;
        RECT 120.420 189.355 134.805 189.455 ;
        RECT 116.420 189.345 117.160 189.355 ;
        RECT 1.100 189.305 19.420 189.325 ;
        RECT 21.010 189.305 21.880 189.325 ;
        RECT 121.190 189.325 134.805 189.355 ;
        RECT 121.190 189.305 122.060 189.325 ;
        RECT 123.650 189.305 134.805 189.325 ;
        RECT 1.100 189.275 18.650 189.305 ;
        RECT 124.420 189.275 134.805 189.305 ;
        RECT 1.100 189.265 18.160 189.275 ;
        RECT 124.910 189.265 134.805 189.275 ;
        RECT 1.100 189.260 17.120 189.265 ;
        RECT 1.100 189.050 2.840 189.260 ;
        RECT 5.170 189.240 17.120 189.260 ;
        RECT 1.020 153.765 2.980 154.180 ;
        RECT 9.985 153.765 10.935 189.240 ;
        RECT 1.020 152.815 10.935 153.765 ;
        RECT 1.020 152.730 2.980 152.815 ;
        RECT 9.985 140.775 10.935 152.815 ;
        RECT 37.745 145.645 38.665 145.975 ;
        RECT 104.405 145.645 105.325 145.975 ;
        RECT 37.730 144.595 38.970 145.015 ;
        RECT 25.920 143.875 38.970 144.595 ;
        RECT 104.100 144.595 105.340 145.015 ;
        RECT 104.100 143.875 117.150 144.595 ;
        RECT 25.920 143.825 38.230 143.875 ;
        RECT 104.840 143.825 117.150 143.875 ;
        RECT 25.920 142.445 26.580 143.825 ;
        RECT 116.490 142.445 117.150 143.825 ;
        RECT 25.910 142.285 26.650 142.445 ;
        RECT 21.230 141.350 22.150 141.680 ;
        RECT 25.920 141.105 26.650 142.285 ;
        RECT 9.985 140.615 17.405 140.775 ;
        RECT 9.985 140.575 18.160 140.615 ;
        RECT 9.985 140.535 18.650 140.575 ;
        RECT 19.300 140.535 21.160 140.555 ;
        RECT 25.910 140.545 26.650 141.105 ;
        RECT 9.985 140.525 21.880 140.535 ;
        RECT 23.900 140.525 26.650 140.545 ;
        RECT 9.985 139.885 26.650 140.525 ;
        RECT 9.985 139.825 22.650 139.885 ;
        RECT 10.000 103.450 10.920 139.825 ;
        RECT 16.360 139.785 22.650 139.825 ;
        RECT 23.580 139.785 26.650 139.885 ;
        RECT 16.360 139.755 21.880 139.785 ;
        RECT 25.910 139.775 26.650 139.785 ;
        RECT 116.420 142.285 117.160 142.445 ;
        RECT 116.420 141.105 117.150 142.285 ;
        RECT 120.920 141.350 121.840 141.680 ;
        RECT 116.420 140.545 117.160 141.105 ;
        RECT 132.315 140.615 134.805 189.265 ;
        RECT 124.910 140.575 134.805 140.615 ;
        RECT 116.420 140.525 119.170 140.545 ;
        RECT 121.910 140.535 123.770 140.555 ;
        RECT 124.420 140.535 134.805 140.575 ;
        RECT 121.190 140.525 134.805 140.535 ;
        RECT 116.420 139.885 134.805 140.525 ;
        RECT 116.420 139.785 119.490 139.885 ;
        RECT 120.420 139.785 134.805 139.885 ;
        RECT 116.420 139.775 117.160 139.785 ;
        RECT 16.360 139.735 19.420 139.755 ;
        RECT 21.010 139.735 21.880 139.755 ;
        RECT 121.190 139.755 134.805 139.785 ;
        RECT 121.190 139.735 122.060 139.755 ;
        RECT 123.650 139.735 134.805 139.755 ;
        RECT 16.360 139.705 18.650 139.735 ;
        RECT 124.420 139.705 134.805 139.735 ;
        RECT 16.360 139.695 18.160 139.705 ;
        RECT 124.910 139.695 134.805 139.705 ;
        RECT 1.070 103.005 3.030 103.420 ;
        RECT 10.000 103.005 10.985 103.450 ;
        RECT 1.070 102.055 10.985 103.005 ;
        RECT 1.070 101.970 3.030 102.055 ;
        RECT 10.000 101.970 10.985 102.055 ;
        RECT 10.000 92.430 10.920 101.970 ;
        RECT 38.405 97.415 39.325 97.745 ;
        RECT 38.390 96.365 39.630 96.785 ;
        RECT 104.405 96.745 105.325 97.075 ;
        RECT 26.580 95.645 39.630 96.365 ;
        RECT 104.100 95.695 105.340 96.115 ;
        RECT 26.580 95.595 38.890 95.645 ;
        RECT 26.580 94.215 27.240 95.595 ;
        RECT 104.100 94.975 117.150 95.695 ;
        RECT 104.840 94.925 117.150 94.975 ;
        RECT 26.570 94.055 27.310 94.215 ;
        RECT 21.890 93.120 22.810 93.450 ;
        RECT 26.580 92.875 27.310 94.055 ;
        RECT 116.490 93.545 117.150 94.925 ;
        RECT 10.000 92.385 18.070 92.430 ;
        RECT 10.000 92.345 18.820 92.385 ;
        RECT 10.000 92.305 19.310 92.345 ;
        RECT 19.960 92.305 21.820 92.325 ;
        RECT 26.570 92.315 27.310 92.875 ;
        RECT 10.000 92.295 22.540 92.305 ;
        RECT 24.560 92.295 27.310 92.315 ;
        RECT 10.000 91.655 27.310 92.295 ;
        RECT 10.000 91.555 23.310 91.655 ;
        RECT 24.240 91.555 27.310 91.655 ;
        RECT 10.000 91.525 22.540 91.555 ;
        RECT 26.570 91.545 27.310 91.555 ;
        RECT 116.420 93.385 117.160 93.545 ;
        RECT 116.420 92.205 117.150 93.385 ;
        RECT 120.920 92.450 121.840 92.780 ;
        RECT 116.420 91.645 117.160 92.205 ;
        RECT 132.315 91.715 134.805 139.695 ;
        RECT 124.910 91.675 134.805 91.715 ;
        RECT 116.420 91.625 119.170 91.645 ;
        RECT 121.910 91.635 123.770 91.655 ;
        RECT 124.420 91.635 134.805 91.675 ;
        RECT 121.190 91.625 134.805 91.635 ;
        RECT 10.000 91.510 20.080 91.525 ;
        RECT 10.015 69.170 10.910 91.510 ;
        RECT 17.020 91.505 20.080 91.510 ;
        RECT 21.670 91.505 22.540 91.525 ;
        RECT 17.020 91.475 19.310 91.505 ;
        RECT 17.020 91.465 18.820 91.475 ;
        RECT 116.420 90.985 134.805 91.625 ;
        RECT 116.420 90.885 119.490 90.985 ;
        RECT 120.420 90.885 134.805 90.985 ;
        RECT 116.420 90.875 117.160 90.885 ;
        RECT 121.190 90.855 134.805 90.885 ;
        RECT 121.190 90.835 122.060 90.855 ;
        RECT 123.650 90.835 134.805 90.855 ;
        RECT 124.420 90.805 134.805 90.835 ;
        RECT 124.910 90.795 134.805 90.805 ;
        RECT 1.030 68.725 2.990 69.140 ;
        RECT 9.995 68.725 10.945 69.170 ;
        RECT 1.030 67.775 10.945 68.725 ;
        RECT 1.030 67.690 2.990 67.775 ;
        RECT 9.995 67.690 10.945 67.775 ;
        RECT 10.015 42.155 10.910 67.690 ;
        RECT 38.075 46.845 38.995 47.175 ;
        RECT 103.745 46.845 104.665 47.175 ;
        RECT 38.060 45.795 39.300 46.215 ;
        RECT 26.250 45.075 39.300 45.795 ;
        RECT 103.440 45.795 104.680 46.215 ;
        RECT 103.440 45.075 116.490 45.795 ;
        RECT 26.250 45.025 38.560 45.075 ;
        RECT 104.180 45.025 116.490 45.075 ;
        RECT 26.250 43.645 26.910 45.025 ;
        RECT 115.830 43.645 116.490 45.025 ;
        RECT 26.240 43.485 26.980 43.645 ;
        RECT 21.560 42.550 22.480 42.880 ;
        RECT 26.250 42.305 26.980 43.485 ;
        RECT 9.840 41.980 11.085 42.155 ;
        RECT 9.840 41.815 17.585 41.980 ;
        RECT 9.840 41.775 18.490 41.815 ;
        RECT 9.840 41.735 18.980 41.775 ;
        RECT 19.630 41.735 21.490 41.755 ;
        RECT 26.240 41.745 26.980 42.305 ;
        RECT 9.840 41.725 22.210 41.735 ;
        RECT 24.230 41.725 26.980 41.745 ;
        RECT 9.840 41.085 26.980 41.725 ;
        RECT 9.840 13.890 11.085 41.085 ;
        RECT 16.690 40.985 22.980 41.085 ;
        RECT 23.910 40.985 26.980 41.085 ;
        RECT 16.690 40.955 22.210 40.985 ;
        RECT 26.240 40.975 26.980 40.985 ;
        RECT 115.760 43.485 116.500 43.645 ;
        RECT 115.760 42.305 116.490 43.485 ;
        RECT 120.260 42.550 121.180 42.880 ;
        RECT 115.760 41.745 116.500 42.305 ;
        RECT 132.315 41.815 134.805 90.795 ;
        RECT 124.250 41.775 134.805 41.815 ;
        RECT 115.760 41.725 118.510 41.745 ;
        RECT 121.250 41.735 123.110 41.755 ;
        RECT 123.760 41.735 134.805 41.775 ;
        RECT 120.530 41.725 134.805 41.735 ;
        RECT 115.760 41.085 134.805 41.725 ;
        RECT 115.760 40.985 118.830 41.085 ;
        RECT 119.760 40.985 134.805 41.085 ;
        RECT 115.760 40.975 116.500 40.985 ;
        RECT 16.690 40.935 19.750 40.955 ;
        RECT 21.340 40.935 22.210 40.955 ;
        RECT 120.530 40.955 134.805 40.985 ;
        RECT 120.530 40.935 121.400 40.955 ;
        RECT 122.990 40.935 134.805 40.955 ;
        RECT 16.690 40.905 18.980 40.935 ;
        RECT 123.760 40.905 134.805 40.935 ;
        RECT 16.690 40.895 18.490 40.905 ;
        RECT 124.250 40.895 134.805 40.905 ;
        RECT 132.315 13.890 134.805 40.895 ;
        RECT 9.220 11.410 134.805 13.890 ;
        RECT 132.315 11.405 134.805 11.410 ;
      LAYER met3 ;
        RECT 37.765 195.205 38.975 195.555 ;
        RECT 104.095 195.205 105.305 195.555 ;
        RECT 37.730 193.445 38.970 194.585 ;
        RECT 104.100 193.445 105.340 194.585 ;
        RECT 20.920 190.910 22.130 191.260 ;
        RECT 120.940 190.910 122.150 191.260 ;
        RECT 1.210 189.265 2.680 190.415 ;
        RECT 18.550 190.040 19.160 190.155 ;
        RECT 18.460 189.330 19.160 190.040 ;
        RECT 18.550 189.225 19.160 189.330 ;
        RECT 21.140 189.265 22.130 190.095 ;
        RECT 120.940 189.265 121.930 190.095 ;
        RECT 123.910 190.040 124.520 190.155 ;
        RECT 123.910 189.330 124.610 190.040 ;
        RECT 123.910 189.225 124.520 189.330 ;
        RECT 1.160 152.835 2.770 153.995 ;
        RECT 37.765 145.635 38.975 145.985 ;
        RECT 104.095 145.635 105.305 145.985 ;
        RECT 37.730 143.875 38.970 145.015 ;
        RECT 104.100 143.875 105.340 145.015 ;
        RECT 20.920 141.340 22.130 141.690 ;
        RECT 120.940 141.340 122.150 141.690 ;
        RECT 18.550 140.470 19.160 140.585 ;
        RECT 18.460 139.760 19.160 140.470 ;
        RECT 18.550 139.655 19.160 139.760 ;
        RECT 21.140 139.695 22.130 140.525 ;
        RECT 120.940 139.695 121.930 140.525 ;
        RECT 123.910 140.470 124.520 140.585 ;
        RECT 123.910 139.760 124.610 140.470 ;
        RECT 123.910 139.655 124.520 139.760 ;
        RECT 1.210 102.075 2.820 103.235 ;
        RECT 38.425 97.405 39.635 97.755 ;
        RECT 38.390 95.645 39.630 96.785 ;
        RECT 104.095 96.735 105.305 97.085 ;
        RECT 104.100 94.975 105.340 96.115 ;
        RECT 21.580 93.110 22.790 93.460 ;
        RECT 120.940 92.440 122.150 92.790 ;
        RECT 19.210 92.240 19.820 92.355 ;
        RECT 19.120 91.530 19.820 92.240 ;
        RECT 19.210 91.425 19.820 91.530 ;
        RECT 21.800 91.465 22.790 92.295 ;
        RECT 120.940 90.795 121.930 91.625 ;
        RECT 123.910 91.570 124.520 91.685 ;
        RECT 123.910 90.860 124.610 91.570 ;
        RECT 123.910 90.755 124.520 90.860 ;
        RECT 1.170 67.795 2.780 68.955 ;
        RECT 38.095 46.835 39.305 47.185 ;
        RECT 103.435 46.835 104.645 47.185 ;
        RECT 38.060 45.075 39.300 46.215 ;
        RECT 103.440 45.075 104.680 46.215 ;
        RECT 21.250 42.540 22.460 42.890 ;
        RECT 120.280 42.540 121.490 42.890 ;
        RECT 18.880 41.670 19.490 41.785 ;
        RECT 18.790 40.960 19.490 41.670 ;
        RECT 18.880 40.855 19.490 40.960 ;
        RECT 21.470 40.895 22.460 41.725 ;
        RECT 120.280 40.895 121.270 41.725 ;
        RECT 123.250 41.670 123.860 41.785 ;
        RECT 123.250 40.960 123.950 41.670 ;
        RECT 123.250 40.855 123.860 40.960 ;
      LAYER met4 ;
        RECT 1.000 103.450 3.000 220.760 ;
        RECT 37.775 194.815 38.975 216.365 ;
        RECT 37.720 194.605 38.975 194.815 ;
        RECT 104.095 194.815 105.295 216.365 ;
        RECT 104.095 194.605 105.350 194.815 ;
        RECT 37.720 193.675 38.970 194.605 ;
        RECT 37.730 193.445 38.970 193.675 ;
        RECT 104.100 193.675 105.350 194.605 ;
        RECT 104.100 193.445 105.340 193.675 ;
        RECT 20.920 170.100 22.120 191.860 ;
        RECT 120.950 170.100 122.150 191.860 ;
        RECT 37.775 145.245 38.975 166.795 ;
        RECT 37.720 145.035 38.975 145.245 ;
        RECT 104.095 145.245 105.295 166.795 ;
        RECT 104.095 145.035 105.350 145.245 ;
        RECT 37.720 144.105 38.970 145.035 ;
        RECT 37.730 143.875 38.970 144.105 ;
        RECT 104.100 144.105 105.350 145.035 ;
        RECT 104.100 143.875 105.340 144.105 ;
        RECT 20.920 120.530 22.120 142.290 ;
        RECT 120.950 120.530 122.150 142.290 ;
        RECT 1.000 101.970 3.050 103.450 ;
        RECT 1.000 69.170 3.000 101.970 ;
        RECT 38.435 97.015 39.635 118.565 ;
        RECT 38.380 96.805 39.635 97.015 ;
        RECT 38.380 95.875 39.630 96.805 ;
        RECT 104.095 96.345 105.295 117.895 ;
        RECT 104.095 96.135 105.350 96.345 ;
        RECT 38.390 95.645 39.630 95.875 ;
        RECT 104.100 95.205 105.350 96.135 ;
        RECT 104.100 94.975 105.340 95.205 ;
        RECT 21.580 72.300 22.780 94.060 ;
        RECT 120.950 71.630 122.150 93.390 ;
        RECT 1.000 67.690 3.010 69.170 ;
        RECT 1.000 5.000 3.000 67.690 ;
        RECT 38.105 46.445 39.305 67.995 ;
        RECT 38.050 46.235 39.305 46.445 ;
        RECT 103.435 46.445 104.635 67.995 ;
        RECT 103.435 46.235 104.690 46.445 ;
        RECT 38.050 45.305 39.300 46.235 ;
        RECT 38.060 45.075 39.300 45.305 ;
        RECT 103.440 45.305 104.690 46.235 ;
        RECT 103.440 45.075 104.680 45.305 ;
        RECT 21.250 21.730 22.450 43.490 ;
        RECT 120.290 21.730 121.490 43.490 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 21.615 194.815 33.085 202.395 ;
        RECT 34.665 201.145 38.695 202.415 ;
        RECT 104.375 201.145 108.405 202.415 ;
        RECT 34.665 197.095 38.695 198.365 ;
        RECT 104.375 197.095 108.405 198.365 ;
        RECT 36.465 195.005 37.525 196.365 ;
        RECT 105.545 195.005 106.605 196.365 ;
        RECT 109.985 194.815 121.455 202.395 ;
        RECT 22.370 190.100 23.430 191.460 ;
        RECT 21.200 188.100 25.230 189.370 ;
      LAYER nwell ;
        RECT 16.715 186.625 18.320 188.035 ;
        RECT 16.715 186.375 18.340 186.625 ;
        RECT 12.460 185.785 13.310 186.305 ;
        RECT 16.690 185.915 18.340 186.375 ;
        RECT 14.820 185.785 18.340 185.915 ;
        RECT 12.460 184.555 18.300 185.785 ;
        RECT 12.460 183.985 13.310 184.555 ;
        RECT 14.820 184.310 18.300 184.555 ;
      LAYER pwell ;
        RECT 21.200 184.050 25.230 185.320 ;
        RECT 26.810 184.070 38.280 191.650 ;
        RECT 104.790 184.070 116.260 191.650 ;
        RECT 119.640 190.100 120.700 191.460 ;
        RECT 117.840 188.100 121.870 189.370 ;
      LAYER nwell ;
        RECT 124.750 186.625 126.355 188.035 ;
        RECT 124.730 186.375 126.355 186.625 ;
        RECT 124.730 185.915 126.380 186.375 ;
        RECT 124.730 185.785 128.250 185.915 ;
        RECT 129.760 185.785 130.610 186.305 ;
      LAYER pwell ;
        RECT 117.840 184.050 121.870 185.320 ;
      LAYER nwell ;
        RECT 124.770 184.555 130.610 185.785 ;
        RECT 124.770 184.310 128.250 184.555 ;
        RECT 129.760 183.985 130.610 184.555 ;
        RECT 12.450 181.685 13.300 182.565 ;
        RECT 16.640 181.805 18.400 181.815 ;
        RECT 14.980 181.685 18.400 181.805 ;
        RECT 12.450 180.505 18.400 181.685 ;
        RECT 12.450 180.245 13.300 180.505 ;
        RECT 14.980 180.210 18.400 180.505 ;
        RECT 124.670 181.805 126.430 181.815 ;
        RECT 124.670 181.685 128.090 181.805 ;
        RECT 129.770 181.685 130.620 182.565 ;
        RECT 124.670 180.505 130.620 181.685 ;
        RECT 124.670 180.210 128.090 180.505 ;
        RECT 129.770 180.245 130.620 180.505 ;
        RECT 14.980 180.200 16.740 180.210 ;
        RECT 126.330 180.200 128.090 180.210 ;
        RECT 16.645 176.665 18.250 178.265 ;
        RECT 16.615 176.505 18.250 176.665 ;
        RECT 124.820 176.665 126.425 178.265 ;
        RECT 124.820 176.505 126.455 176.665 ;
        RECT 16.615 175.385 18.220 176.505 ;
        RECT 16.610 175.105 18.220 175.385 ;
        RECT 124.850 175.385 126.455 176.505 ;
        RECT 124.850 175.105 126.460 175.385 ;
        RECT 16.610 174.765 18.280 175.105 ;
        RECT 124.790 174.765 126.460 175.105 ;
        RECT 16.610 173.905 18.290 174.765 ;
        RECT 15.500 173.115 18.290 173.905 ;
        RECT 124.780 173.905 126.460 174.765 ;
        RECT 124.780 173.115 127.570 173.905 ;
        RECT 15.500 173.065 18.260 173.115 ;
        RECT 124.810 173.065 127.570 173.115 ;
        RECT 15.500 173.055 17.820 173.065 ;
        RECT 125.250 173.055 127.570 173.065 ;
      LAYER pwell ;
        RECT 21.615 145.245 33.085 152.825 ;
        RECT 34.665 151.575 38.695 152.845 ;
        RECT 104.375 151.575 108.405 152.845 ;
        RECT 34.665 147.525 38.695 148.795 ;
        RECT 104.375 147.525 108.405 148.795 ;
        RECT 36.465 145.435 37.525 146.795 ;
        RECT 105.545 145.435 106.605 146.795 ;
        RECT 109.985 145.245 121.455 152.825 ;
        RECT 22.370 140.530 23.430 141.890 ;
        RECT 21.200 138.530 25.230 139.800 ;
      LAYER nwell ;
        RECT 16.715 137.055 18.320 138.465 ;
        RECT 16.715 136.805 18.340 137.055 ;
        RECT 12.460 136.215 13.310 136.735 ;
        RECT 16.690 136.345 18.340 136.805 ;
        RECT 14.820 136.215 18.340 136.345 ;
        RECT 12.460 134.985 18.300 136.215 ;
        RECT 12.460 134.415 13.310 134.985 ;
        RECT 14.820 134.740 18.300 134.985 ;
      LAYER pwell ;
        RECT 21.200 134.480 25.230 135.750 ;
        RECT 26.810 134.500 38.280 142.080 ;
        RECT 104.790 134.500 116.260 142.080 ;
        RECT 119.640 140.530 120.700 141.890 ;
        RECT 117.840 138.530 121.870 139.800 ;
      LAYER nwell ;
        RECT 124.750 137.055 126.355 138.465 ;
        RECT 124.730 136.805 126.355 137.055 ;
        RECT 124.730 136.345 126.380 136.805 ;
        RECT 124.730 136.215 128.250 136.345 ;
        RECT 129.760 136.215 130.610 136.735 ;
      LAYER pwell ;
        RECT 117.840 134.480 121.870 135.750 ;
      LAYER nwell ;
        RECT 124.770 134.985 130.610 136.215 ;
        RECT 124.770 134.740 128.250 134.985 ;
        RECT 129.760 134.415 130.610 134.985 ;
        RECT 12.450 132.115 13.300 132.995 ;
        RECT 16.640 132.235 18.400 132.245 ;
        RECT 14.980 132.115 18.400 132.235 ;
        RECT 12.450 130.935 18.400 132.115 ;
        RECT 12.450 130.675 13.300 130.935 ;
        RECT 14.980 130.640 18.400 130.935 ;
        RECT 124.670 132.235 126.430 132.245 ;
        RECT 124.670 132.115 128.090 132.235 ;
        RECT 129.770 132.115 130.620 132.995 ;
        RECT 124.670 130.935 130.620 132.115 ;
        RECT 124.670 130.640 128.090 130.935 ;
        RECT 129.770 130.675 130.620 130.935 ;
        RECT 14.980 130.630 16.740 130.640 ;
        RECT 126.330 130.630 128.090 130.640 ;
        RECT 16.645 127.095 18.250 128.695 ;
        RECT 16.615 126.935 18.250 127.095 ;
        RECT 124.820 127.095 126.425 128.695 ;
        RECT 124.820 126.935 126.455 127.095 ;
        RECT 16.615 125.815 18.220 126.935 ;
        RECT 16.610 125.535 18.220 125.815 ;
        RECT 124.850 125.815 126.455 126.935 ;
        RECT 124.850 125.535 126.460 125.815 ;
        RECT 16.610 125.195 18.280 125.535 ;
        RECT 124.790 125.195 126.460 125.535 ;
        RECT 16.610 124.335 18.290 125.195 ;
        RECT 15.500 123.545 18.290 124.335 ;
        RECT 124.780 124.335 126.460 125.195 ;
        RECT 124.780 123.545 127.570 124.335 ;
        RECT 15.500 123.495 18.260 123.545 ;
        RECT 124.810 123.495 127.570 123.545 ;
        RECT 15.500 123.485 17.820 123.495 ;
        RECT 125.250 123.485 127.570 123.495 ;
      LAYER pwell ;
        RECT 22.275 97.015 33.745 104.595 ;
        RECT 35.325 103.345 39.355 104.615 ;
        RECT 104.375 102.675 108.405 103.945 ;
        RECT 35.325 99.295 39.355 100.565 ;
        RECT 104.375 98.625 108.405 99.895 ;
        RECT 37.125 97.205 38.185 98.565 ;
        RECT 105.545 96.535 106.605 97.895 ;
        RECT 109.985 96.345 121.455 103.925 ;
        RECT 23.030 92.300 24.090 93.660 ;
        RECT 21.860 90.300 25.890 91.570 ;
      LAYER nwell ;
        RECT 17.375 88.825 18.980 90.235 ;
        RECT 17.375 88.575 19.000 88.825 ;
        RECT 13.120 87.985 13.970 88.505 ;
        RECT 17.350 88.115 19.000 88.575 ;
        RECT 15.480 87.985 19.000 88.115 ;
        RECT 13.120 86.755 18.960 87.985 ;
        RECT 13.120 86.185 13.970 86.755 ;
        RECT 15.480 86.510 18.960 86.755 ;
      LAYER pwell ;
        RECT 21.860 86.250 25.890 87.520 ;
        RECT 27.470 86.270 38.940 93.850 ;
        RECT 104.790 85.600 116.260 93.180 ;
        RECT 119.640 91.630 120.700 92.990 ;
        RECT 117.840 89.630 121.870 90.900 ;
      LAYER nwell ;
        RECT 124.750 88.155 126.355 89.565 ;
        RECT 124.730 87.905 126.355 88.155 ;
        RECT 124.730 87.445 126.380 87.905 ;
        RECT 124.730 87.315 128.250 87.445 ;
        RECT 129.760 87.315 130.610 87.835 ;
      LAYER pwell ;
        RECT 117.840 85.580 121.870 86.850 ;
      LAYER nwell ;
        RECT 124.770 86.085 130.610 87.315 ;
        RECT 124.770 85.840 128.250 86.085 ;
        RECT 129.760 85.515 130.610 86.085 ;
        RECT 13.110 83.885 13.960 84.765 ;
        RECT 17.300 84.005 19.060 84.015 ;
        RECT 15.640 83.885 19.060 84.005 ;
        RECT 13.110 82.705 19.060 83.885 ;
        RECT 13.110 82.445 13.960 82.705 ;
        RECT 15.640 82.410 19.060 82.705 ;
        RECT 124.670 83.335 126.430 83.345 ;
        RECT 124.670 83.215 128.090 83.335 ;
        RECT 129.770 83.215 130.620 84.095 ;
        RECT 15.640 82.400 17.400 82.410 ;
        RECT 124.670 82.035 130.620 83.215 ;
        RECT 124.670 81.740 128.090 82.035 ;
        RECT 129.770 81.775 130.620 82.035 ;
        RECT 126.330 81.730 128.090 81.740 ;
        RECT 17.305 78.865 18.910 80.465 ;
        RECT 17.275 78.705 18.910 78.865 ;
        RECT 17.275 77.585 18.880 78.705 ;
        RECT 124.820 78.195 126.425 79.795 ;
        RECT 124.820 78.035 126.455 78.195 ;
        RECT 17.270 77.305 18.880 77.585 ;
        RECT 17.270 76.965 18.940 77.305 ;
        RECT 17.270 76.105 18.950 76.965 ;
        RECT 124.850 76.915 126.455 78.035 ;
        RECT 124.850 76.635 126.460 76.915 ;
        RECT 124.790 76.295 126.460 76.635 ;
        RECT 16.160 75.315 18.950 76.105 ;
        RECT 124.780 75.435 126.460 76.295 ;
        RECT 16.160 75.265 18.920 75.315 ;
        RECT 16.160 75.255 18.480 75.265 ;
        RECT 124.780 74.645 127.570 75.435 ;
        RECT 124.810 74.595 127.570 74.645 ;
        RECT 125.250 74.585 127.570 74.595 ;
      LAYER pwell ;
        RECT 21.945 46.445 33.415 54.025 ;
        RECT 34.995 52.775 39.025 54.045 ;
        RECT 103.715 52.775 107.745 54.045 ;
        RECT 34.995 48.725 39.025 49.995 ;
        RECT 103.715 48.725 107.745 49.995 ;
        RECT 36.795 46.635 37.855 47.995 ;
        RECT 104.885 46.635 105.945 47.995 ;
        RECT 109.325 46.445 120.795 54.025 ;
        RECT 22.700 41.730 23.760 43.090 ;
        RECT 21.530 39.730 25.560 41.000 ;
      LAYER nwell ;
        RECT 17.045 38.255 18.650 39.665 ;
        RECT 17.045 38.005 18.670 38.255 ;
        RECT 12.790 37.415 13.640 37.935 ;
        RECT 17.020 37.545 18.670 38.005 ;
        RECT 15.150 37.415 18.670 37.545 ;
        RECT 12.790 36.185 18.630 37.415 ;
        RECT 12.790 35.615 13.640 36.185 ;
        RECT 15.150 35.940 18.630 36.185 ;
      LAYER pwell ;
        RECT 21.530 35.680 25.560 36.950 ;
        RECT 27.140 35.700 38.610 43.280 ;
        RECT 104.130 35.700 115.600 43.280 ;
        RECT 118.980 41.730 120.040 43.090 ;
        RECT 117.180 39.730 121.210 41.000 ;
      LAYER nwell ;
        RECT 124.090 38.255 125.695 39.665 ;
        RECT 124.070 38.005 125.695 38.255 ;
        RECT 124.070 37.545 125.720 38.005 ;
        RECT 124.070 37.415 127.590 37.545 ;
        RECT 129.100 37.415 129.950 37.935 ;
      LAYER pwell ;
        RECT 117.180 35.680 121.210 36.950 ;
      LAYER nwell ;
        RECT 124.110 36.185 129.950 37.415 ;
        RECT 124.110 35.940 127.590 36.185 ;
        RECT 129.100 35.615 129.950 36.185 ;
        RECT 12.780 33.315 13.630 34.195 ;
        RECT 16.970 33.435 18.730 33.445 ;
        RECT 15.310 33.315 18.730 33.435 ;
        RECT 12.780 32.135 18.730 33.315 ;
        RECT 12.780 31.875 13.630 32.135 ;
        RECT 15.310 31.840 18.730 32.135 ;
        RECT 124.010 33.435 125.770 33.445 ;
        RECT 124.010 33.315 127.430 33.435 ;
        RECT 129.110 33.315 129.960 34.195 ;
        RECT 124.010 32.135 129.960 33.315 ;
        RECT 124.010 31.840 127.430 32.135 ;
        RECT 129.110 31.875 129.960 32.135 ;
        RECT 15.310 31.830 17.070 31.840 ;
        RECT 125.670 31.830 127.430 31.840 ;
        RECT 16.975 28.295 18.580 29.895 ;
        RECT 16.945 28.135 18.580 28.295 ;
        RECT 124.160 28.295 125.765 29.895 ;
        RECT 124.160 28.135 125.795 28.295 ;
        RECT 16.945 27.015 18.550 28.135 ;
        RECT 16.940 26.735 18.550 27.015 ;
        RECT 124.190 27.015 125.795 28.135 ;
        RECT 124.190 26.735 125.800 27.015 ;
        RECT 16.940 26.395 18.610 26.735 ;
        RECT 124.130 26.395 125.800 26.735 ;
        RECT 16.940 25.535 18.620 26.395 ;
        RECT 15.830 24.745 18.620 25.535 ;
        RECT 124.120 25.535 125.800 26.395 ;
        RECT 124.120 24.745 126.910 25.535 ;
        RECT 15.830 24.695 18.590 24.745 ;
        RECT 124.150 24.695 126.910 24.745 ;
        RECT 15.830 24.685 18.150 24.695 ;
        RECT 124.590 24.685 126.910 24.695 ;
      LAYER li1 ;
        RECT 21.855 201.985 32.845 202.155 ;
        RECT 21.855 195.225 22.025 201.985 ;
        RECT 32.675 195.225 32.845 201.985 ;
        RECT 35.205 201.585 35.375 202.115 ;
        RECT 36.555 201.525 37.595 201.865 ;
        RECT 105.475 201.525 106.515 201.865 ;
        RECT 107.695 201.585 107.865 202.115 ;
        RECT 110.225 201.985 121.215 202.155 ;
        RECT 35.205 197.395 35.375 197.925 ;
        RECT 36.555 197.645 37.595 197.985 ;
        RECT 105.475 197.645 106.515 197.985 ;
        RECT 107.695 197.395 107.865 197.925 ;
        RECT 21.855 195.055 32.845 195.225 ;
        RECT 36.685 195.115 37.025 195.785 ;
        RECT 106.045 195.115 106.385 195.785 ;
        RECT 110.225 195.225 110.395 201.985 ;
        RECT 121.045 195.225 121.215 201.985 ;
        RECT 110.225 195.055 121.215 195.225 ;
        RECT 22.870 190.680 23.210 191.350 ;
        RECT 27.050 191.240 38.040 191.410 ;
        RECT 22.300 188.480 23.340 188.820 ;
        RECT 24.520 188.540 24.690 189.070 ;
        RECT 15.325 187.750 15.495 187.845 ;
        RECT 15.325 187.480 16.305 187.750 ;
        RECT 15.325 186.810 15.495 187.480 ;
        RECT 15.325 186.570 16.305 186.810 ;
        RECT 15.325 186.465 15.495 186.570 ;
        RECT 12.655 185.950 12.840 186.120 ;
        RECT 12.655 185.435 12.825 185.950 ;
        RECT 14.380 185.435 14.900 185.465 ;
        RECT 12.655 184.875 14.900 185.435 ;
        RECT 12.640 184.845 14.900 184.875 ;
        RECT 12.640 184.835 14.750 184.845 ;
        RECT 12.640 181.625 12.850 184.835 ;
        RECT 22.300 184.600 23.340 184.940 ;
        RECT 24.520 184.350 24.690 184.880 ;
        RECT 27.050 184.480 27.220 191.240 ;
        RECT 28.510 185.340 28.680 190.380 ;
        RECT 30.090 185.340 30.260 190.380 ;
        RECT 31.670 185.340 31.840 190.380 ;
        RECT 33.250 185.340 33.420 190.380 ;
        RECT 34.830 185.340 35.000 190.380 ;
        RECT 36.410 185.340 36.580 190.380 ;
        RECT 37.870 184.480 38.040 191.240 ;
        RECT 27.050 184.310 38.040 184.480 ;
        RECT 105.030 191.240 116.020 191.410 ;
        RECT 105.030 184.480 105.200 191.240 ;
        RECT 106.490 185.340 106.660 190.380 ;
        RECT 108.070 185.340 108.240 190.380 ;
        RECT 109.650 185.340 109.820 190.380 ;
        RECT 111.230 185.340 111.400 190.380 ;
        RECT 112.810 185.340 112.980 190.380 ;
        RECT 114.390 185.340 114.560 190.380 ;
        RECT 115.850 184.480 116.020 191.240 ;
        RECT 119.860 190.680 120.200 191.350 ;
        RECT 118.380 188.540 118.550 189.070 ;
        RECT 119.730 188.480 120.770 188.820 ;
        RECT 127.575 187.750 127.745 187.845 ;
        RECT 126.765 187.480 127.745 187.750 ;
        RECT 127.575 186.810 127.745 187.480 ;
        RECT 126.765 186.570 127.745 186.810 ;
        RECT 127.575 186.465 127.745 186.570 ;
        RECT 130.230 185.950 130.415 186.120 ;
        RECT 128.170 185.435 128.690 185.465 ;
        RECT 130.245 185.435 130.415 185.950 ;
        RECT 105.030 184.310 116.020 184.480 ;
        RECT 118.380 184.350 118.550 184.880 ;
        RECT 119.730 184.600 120.770 184.940 ;
        RECT 128.170 184.875 130.415 185.435 ;
        RECT 128.170 184.845 130.430 184.875 ;
        RECT 128.320 184.835 130.430 184.845 ;
        RECT 15.840 183.090 16.070 183.910 ;
        RECT 17.560 183.090 17.790 183.910 ;
        RECT 125.280 183.090 125.510 183.910 ;
        RECT 127.000 183.090 127.230 183.910 ;
        RECT 15.010 182.920 16.390 183.090 ;
        RECT 16.730 182.920 18.110 183.090 ;
        RECT 124.960 182.920 126.340 183.090 ;
        RECT 126.680 182.920 128.060 183.090 ;
        RECT 12.645 180.600 12.815 181.625 ;
        RECT 12.645 180.430 12.830 180.600 ;
        RECT 16.000 178.980 16.230 179.800 ;
        RECT 17.660 178.990 17.890 179.810 ;
        RECT 15.170 178.810 16.550 178.980 ;
        RECT 16.830 178.820 18.210 178.990 ;
        RECT 15.255 177.980 15.425 178.075 ;
        RECT 15.255 177.710 16.235 177.980 ;
        RECT 15.255 177.040 15.425 177.710 ;
        RECT 15.255 176.800 16.235 177.040 ;
        RECT 15.255 176.695 15.425 176.800 ;
        RECT 15.225 175.645 15.395 176.475 ;
        RECT 15.225 175.415 16.215 175.645 ;
        RECT 15.225 175.405 15.395 175.415 ;
        RECT 15.210 175.095 15.395 175.405 ;
        RECT 15.210 173.705 15.390 175.095 ;
        RECT 17.460 173.710 17.790 173.715 ;
        RECT 15.685 173.705 17.790 173.710 ;
        RECT 15.210 173.540 17.790 173.705 ;
        RECT 15.210 173.525 15.855 173.540 ;
        RECT 17.460 173.535 17.790 173.540 ;
        RECT 17.465 173.525 17.635 173.535 ;
        RECT 15.210 173.495 15.840 173.525 ;
        RECT 15.220 173.485 15.840 173.495 ;
        RECT 23.620 171.815 23.790 181.855 ;
        RECT 25.200 171.815 25.370 181.855 ;
        RECT 26.780 171.815 26.950 181.855 ;
        RECT 28.360 171.815 28.530 181.855 ;
        RECT 29.940 171.815 30.110 181.855 ;
        RECT 31.520 171.815 31.690 181.855 ;
        RECT 33.100 171.815 33.270 181.855 ;
        RECT 34.680 171.815 34.850 181.855 ;
        RECT 36.260 171.815 36.430 181.855 ;
        RECT 106.640 171.815 106.810 181.855 ;
        RECT 108.220 171.815 108.390 181.855 ;
        RECT 109.800 171.815 109.970 181.855 ;
        RECT 111.380 171.815 111.550 181.855 ;
        RECT 112.960 171.815 113.130 181.855 ;
        RECT 114.540 171.815 114.710 181.855 ;
        RECT 116.120 171.815 116.290 181.855 ;
        RECT 117.700 171.815 117.870 181.855 ;
        RECT 119.280 171.815 119.450 181.855 ;
        RECT 130.220 181.625 130.430 184.835 ;
        RECT 130.255 180.600 130.425 181.625 ;
        RECT 130.240 180.430 130.425 180.600 ;
        RECT 125.180 178.990 125.410 179.810 ;
        RECT 124.860 178.820 126.240 178.990 ;
        RECT 126.840 178.980 127.070 179.800 ;
        RECT 126.520 178.810 127.900 178.980 ;
        RECT 127.645 177.980 127.815 178.075 ;
        RECT 126.835 177.710 127.815 177.980 ;
        RECT 127.645 177.040 127.815 177.710 ;
        RECT 126.835 176.800 127.815 177.040 ;
        RECT 127.645 176.695 127.815 176.800 ;
        RECT 127.675 175.645 127.845 176.475 ;
        RECT 126.855 175.415 127.845 175.645 ;
        RECT 127.675 175.405 127.845 175.415 ;
        RECT 127.675 175.095 127.860 175.405 ;
        RECT 125.280 173.710 125.610 173.715 ;
        RECT 125.280 173.705 127.385 173.710 ;
        RECT 127.680 173.705 127.860 175.095 ;
        RECT 125.280 173.540 127.860 173.705 ;
        RECT 125.280 173.535 125.610 173.540 ;
        RECT 125.435 173.525 125.605 173.535 ;
        RECT 127.215 173.525 127.860 173.540 ;
        RECT 127.230 173.495 127.860 173.525 ;
        RECT 127.230 173.485 127.850 173.495 ;
        RECT 21.855 152.415 32.845 152.585 ;
        RECT 21.855 145.655 22.025 152.415 ;
        RECT 32.675 145.655 32.845 152.415 ;
        RECT 35.205 152.015 35.375 152.545 ;
        RECT 36.555 151.955 37.595 152.295 ;
        RECT 105.475 151.955 106.515 152.295 ;
        RECT 107.695 152.015 107.865 152.545 ;
        RECT 110.225 152.415 121.215 152.585 ;
        RECT 35.205 147.825 35.375 148.355 ;
        RECT 36.555 148.075 37.595 148.415 ;
        RECT 105.475 148.075 106.515 148.415 ;
        RECT 107.695 147.825 107.865 148.355 ;
        RECT 21.855 145.485 32.845 145.655 ;
        RECT 36.685 145.545 37.025 146.215 ;
        RECT 106.045 145.545 106.385 146.215 ;
        RECT 110.225 145.655 110.395 152.415 ;
        RECT 121.045 145.655 121.215 152.415 ;
        RECT 110.225 145.485 121.215 145.655 ;
        RECT 22.870 141.110 23.210 141.780 ;
        RECT 27.050 141.670 38.040 141.840 ;
        RECT 22.300 138.910 23.340 139.250 ;
        RECT 24.520 138.970 24.690 139.500 ;
        RECT 15.325 138.180 15.495 138.275 ;
        RECT 15.325 137.910 16.305 138.180 ;
        RECT 15.325 137.240 15.495 137.910 ;
        RECT 15.325 137.000 16.305 137.240 ;
        RECT 15.325 136.895 15.495 137.000 ;
        RECT 12.655 136.380 12.840 136.550 ;
        RECT 12.655 135.865 12.825 136.380 ;
        RECT 14.380 135.865 14.900 135.895 ;
        RECT 12.655 135.305 14.900 135.865 ;
        RECT 12.640 135.275 14.900 135.305 ;
        RECT 12.640 135.265 14.750 135.275 ;
        RECT 12.640 132.055 12.850 135.265 ;
        RECT 22.300 135.030 23.340 135.370 ;
        RECT 24.520 134.780 24.690 135.310 ;
        RECT 27.050 134.910 27.220 141.670 ;
        RECT 28.510 135.770 28.680 140.810 ;
        RECT 30.090 135.770 30.260 140.810 ;
        RECT 31.670 135.770 31.840 140.810 ;
        RECT 33.250 135.770 33.420 140.810 ;
        RECT 34.830 135.770 35.000 140.810 ;
        RECT 36.410 135.770 36.580 140.810 ;
        RECT 37.870 134.910 38.040 141.670 ;
        RECT 27.050 134.740 38.040 134.910 ;
        RECT 105.030 141.670 116.020 141.840 ;
        RECT 105.030 134.910 105.200 141.670 ;
        RECT 106.490 135.770 106.660 140.810 ;
        RECT 108.070 135.770 108.240 140.810 ;
        RECT 109.650 135.770 109.820 140.810 ;
        RECT 111.230 135.770 111.400 140.810 ;
        RECT 112.810 135.770 112.980 140.810 ;
        RECT 114.390 135.770 114.560 140.810 ;
        RECT 115.850 134.910 116.020 141.670 ;
        RECT 119.860 141.110 120.200 141.780 ;
        RECT 118.380 138.970 118.550 139.500 ;
        RECT 119.730 138.910 120.770 139.250 ;
        RECT 127.575 138.180 127.745 138.275 ;
        RECT 126.765 137.910 127.745 138.180 ;
        RECT 127.575 137.240 127.745 137.910 ;
        RECT 126.765 137.000 127.745 137.240 ;
        RECT 127.575 136.895 127.745 137.000 ;
        RECT 130.230 136.380 130.415 136.550 ;
        RECT 128.170 135.865 128.690 135.895 ;
        RECT 130.245 135.865 130.415 136.380 ;
        RECT 105.030 134.740 116.020 134.910 ;
        RECT 118.380 134.780 118.550 135.310 ;
        RECT 119.730 135.030 120.770 135.370 ;
        RECT 128.170 135.305 130.415 135.865 ;
        RECT 128.170 135.275 130.430 135.305 ;
        RECT 128.320 135.265 130.430 135.275 ;
        RECT 15.840 133.520 16.070 134.340 ;
        RECT 17.560 133.520 17.790 134.340 ;
        RECT 125.280 133.520 125.510 134.340 ;
        RECT 127.000 133.520 127.230 134.340 ;
        RECT 15.010 133.350 16.390 133.520 ;
        RECT 16.730 133.350 18.110 133.520 ;
        RECT 124.960 133.350 126.340 133.520 ;
        RECT 126.680 133.350 128.060 133.520 ;
        RECT 12.645 131.030 12.815 132.055 ;
        RECT 12.645 130.860 12.830 131.030 ;
        RECT 16.000 129.410 16.230 130.230 ;
        RECT 17.660 129.420 17.890 130.240 ;
        RECT 15.170 129.240 16.550 129.410 ;
        RECT 16.830 129.250 18.210 129.420 ;
        RECT 15.255 128.410 15.425 128.505 ;
        RECT 15.255 128.140 16.235 128.410 ;
        RECT 15.255 127.470 15.425 128.140 ;
        RECT 15.255 127.230 16.235 127.470 ;
        RECT 15.255 127.125 15.425 127.230 ;
        RECT 15.225 126.075 15.395 126.905 ;
        RECT 15.225 125.845 16.215 126.075 ;
        RECT 15.225 125.835 15.395 125.845 ;
        RECT 15.210 125.525 15.395 125.835 ;
        RECT 15.210 124.135 15.390 125.525 ;
        RECT 17.460 124.140 17.790 124.145 ;
        RECT 15.685 124.135 17.790 124.140 ;
        RECT 15.210 123.970 17.790 124.135 ;
        RECT 15.210 123.955 15.855 123.970 ;
        RECT 17.460 123.965 17.790 123.970 ;
        RECT 17.465 123.955 17.635 123.965 ;
        RECT 15.210 123.925 15.840 123.955 ;
        RECT 15.220 123.915 15.840 123.925 ;
        RECT 23.620 122.245 23.790 132.285 ;
        RECT 25.200 122.245 25.370 132.285 ;
        RECT 26.780 122.245 26.950 132.285 ;
        RECT 28.360 122.245 28.530 132.285 ;
        RECT 29.940 122.245 30.110 132.285 ;
        RECT 31.520 122.245 31.690 132.285 ;
        RECT 33.100 122.245 33.270 132.285 ;
        RECT 34.680 122.245 34.850 132.285 ;
        RECT 36.260 122.245 36.430 132.285 ;
        RECT 106.640 122.245 106.810 132.285 ;
        RECT 108.220 122.245 108.390 132.285 ;
        RECT 109.800 122.245 109.970 132.285 ;
        RECT 111.380 122.245 111.550 132.285 ;
        RECT 112.960 122.245 113.130 132.285 ;
        RECT 114.540 122.245 114.710 132.285 ;
        RECT 116.120 122.245 116.290 132.285 ;
        RECT 117.700 122.245 117.870 132.285 ;
        RECT 119.280 122.245 119.450 132.285 ;
        RECT 130.220 132.055 130.430 135.265 ;
        RECT 130.255 131.030 130.425 132.055 ;
        RECT 130.240 130.860 130.425 131.030 ;
        RECT 125.180 129.420 125.410 130.240 ;
        RECT 124.860 129.250 126.240 129.420 ;
        RECT 126.840 129.410 127.070 130.230 ;
        RECT 126.520 129.240 127.900 129.410 ;
        RECT 127.645 128.410 127.815 128.505 ;
        RECT 126.835 128.140 127.815 128.410 ;
        RECT 127.645 127.470 127.815 128.140 ;
        RECT 126.835 127.230 127.815 127.470 ;
        RECT 127.645 127.125 127.815 127.230 ;
        RECT 127.675 126.075 127.845 126.905 ;
        RECT 126.855 125.845 127.845 126.075 ;
        RECT 127.675 125.835 127.845 125.845 ;
        RECT 127.675 125.525 127.860 125.835 ;
        RECT 125.280 124.140 125.610 124.145 ;
        RECT 125.280 124.135 127.385 124.140 ;
        RECT 127.680 124.135 127.860 125.525 ;
        RECT 125.280 123.970 127.860 124.135 ;
        RECT 125.280 123.965 125.610 123.970 ;
        RECT 125.435 123.955 125.605 123.965 ;
        RECT 127.215 123.955 127.860 123.970 ;
        RECT 127.230 123.925 127.860 123.955 ;
        RECT 127.230 123.915 127.850 123.925 ;
        RECT 22.515 104.185 33.505 104.355 ;
        RECT 22.515 97.425 22.685 104.185 ;
        RECT 33.335 97.425 33.505 104.185 ;
        RECT 35.865 103.785 36.035 104.315 ;
        RECT 37.215 103.725 38.255 104.065 ;
        RECT 105.475 103.055 106.515 103.395 ;
        RECT 107.695 103.115 107.865 103.645 ;
        RECT 110.225 103.515 121.215 103.685 ;
        RECT 35.865 99.595 36.035 100.125 ;
        RECT 37.215 99.845 38.255 100.185 ;
        RECT 105.475 99.175 106.515 99.515 ;
        RECT 107.695 98.925 107.865 99.455 ;
        RECT 22.515 97.255 33.505 97.425 ;
        RECT 37.345 97.315 37.685 97.985 ;
        RECT 106.045 96.645 106.385 97.315 ;
        RECT 110.225 96.755 110.395 103.515 ;
        RECT 121.045 96.755 121.215 103.515 ;
        RECT 110.225 96.585 121.215 96.755 ;
        RECT 23.530 92.880 23.870 93.550 ;
        RECT 27.710 93.440 38.700 93.610 ;
        RECT 22.960 90.680 24.000 91.020 ;
        RECT 25.180 90.740 25.350 91.270 ;
        RECT 15.985 89.950 16.155 90.045 ;
        RECT 15.985 89.680 16.965 89.950 ;
        RECT 15.985 89.010 16.155 89.680 ;
        RECT 15.985 88.770 16.965 89.010 ;
        RECT 15.985 88.665 16.155 88.770 ;
        RECT 13.315 88.150 13.500 88.320 ;
        RECT 13.315 87.635 13.485 88.150 ;
        RECT 15.040 87.635 15.560 87.665 ;
        RECT 13.315 87.075 15.560 87.635 ;
        RECT 13.300 87.045 15.560 87.075 ;
        RECT 13.300 87.035 15.410 87.045 ;
        RECT 13.300 83.825 13.510 87.035 ;
        RECT 22.960 86.800 24.000 87.140 ;
        RECT 25.180 86.550 25.350 87.080 ;
        RECT 27.710 86.680 27.880 93.440 ;
        RECT 29.170 87.540 29.340 92.580 ;
        RECT 30.750 87.540 30.920 92.580 ;
        RECT 32.330 87.540 32.500 92.580 ;
        RECT 33.910 87.540 34.080 92.580 ;
        RECT 35.490 87.540 35.660 92.580 ;
        RECT 37.070 87.540 37.240 92.580 ;
        RECT 38.530 86.680 38.700 93.440 ;
        RECT 27.710 86.510 38.700 86.680 ;
        RECT 105.030 92.770 116.020 92.940 ;
        RECT 16.500 85.290 16.730 86.110 ;
        RECT 18.220 85.290 18.450 86.110 ;
        RECT 105.030 86.010 105.200 92.770 ;
        RECT 106.490 86.870 106.660 91.910 ;
        RECT 108.070 86.870 108.240 91.910 ;
        RECT 109.650 86.870 109.820 91.910 ;
        RECT 111.230 86.870 111.400 91.910 ;
        RECT 112.810 86.870 112.980 91.910 ;
        RECT 114.390 86.870 114.560 91.910 ;
        RECT 115.850 86.010 116.020 92.770 ;
        RECT 119.860 92.210 120.200 92.880 ;
        RECT 118.380 90.070 118.550 90.600 ;
        RECT 119.730 90.010 120.770 90.350 ;
        RECT 127.575 89.280 127.745 89.375 ;
        RECT 126.765 89.010 127.745 89.280 ;
        RECT 127.575 88.340 127.745 89.010 ;
        RECT 126.765 88.100 127.745 88.340 ;
        RECT 127.575 87.995 127.745 88.100 ;
        RECT 130.230 87.480 130.415 87.650 ;
        RECT 128.170 86.965 128.690 86.995 ;
        RECT 130.245 86.965 130.415 87.480 ;
        RECT 105.030 85.840 116.020 86.010 ;
        RECT 118.380 85.880 118.550 86.410 ;
        RECT 119.730 86.130 120.770 86.470 ;
        RECT 128.170 86.405 130.415 86.965 ;
        RECT 128.170 86.375 130.430 86.405 ;
        RECT 128.320 86.365 130.430 86.375 ;
        RECT 15.670 85.120 17.050 85.290 ;
        RECT 17.390 85.120 18.770 85.290 ;
        RECT 125.280 84.620 125.510 85.440 ;
        RECT 127.000 84.620 127.230 85.440 ;
        RECT 124.960 84.450 126.340 84.620 ;
        RECT 126.680 84.450 128.060 84.620 ;
        RECT 13.305 82.800 13.475 83.825 ;
        RECT 13.305 82.630 13.490 82.800 ;
        RECT 16.660 81.180 16.890 82.000 ;
        RECT 18.320 81.190 18.550 82.010 ;
        RECT 15.830 81.010 17.210 81.180 ;
        RECT 17.490 81.020 18.870 81.190 ;
        RECT 15.915 80.180 16.085 80.275 ;
        RECT 15.915 79.910 16.895 80.180 ;
        RECT 15.915 79.240 16.085 79.910 ;
        RECT 15.915 79.000 16.895 79.240 ;
        RECT 15.915 78.895 16.085 79.000 ;
        RECT 15.885 77.845 16.055 78.675 ;
        RECT 15.885 77.615 16.875 77.845 ;
        RECT 15.885 77.605 16.055 77.615 ;
        RECT 15.870 77.295 16.055 77.605 ;
        RECT 15.870 75.905 16.050 77.295 ;
        RECT 18.120 75.910 18.450 75.915 ;
        RECT 16.345 75.905 18.450 75.910 ;
        RECT 15.870 75.740 18.450 75.905 ;
        RECT 15.870 75.725 16.515 75.740 ;
        RECT 18.120 75.735 18.450 75.740 ;
        RECT 18.125 75.725 18.295 75.735 ;
        RECT 15.870 75.695 16.500 75.725 ;
        RECT 15.880 75.685 16.500 75.695 ;
        RECT 24.280 74.015 24.450 84.055 ;
        RECT 25.860 74.015 26.030 84.055 ;
        RECT 27.440 74.015 27.610 84.055 ;
        RECT 29.020 74.015 29.190 84.055 ;
        RECT 30.600 74.015 30.770 84.055 ;
        RECT 32.180 74.015 32.350 84.055 ;
        RECT 33.760 74.015 33.930 84.055 ;
        RECT 35.340 74.015 35.510 84.055 ;
        RECT 36.920 74.015 37.090 84.055 ;
        RECT 106.640 73.345 106.810 83.385 ;
        RECT 108.220 73.345 108.390 83.385 ;
        RECT 109.800 73.345 109.970 83.385 ;
        RECT 111.380 73.345 111.550 83.385 ;
        RECT 112.960 73.345 113.130 83.385 ;
        RECT 114.540 73.345 114.710 83.385 ;
        RECT 116.120 73.345 116.290 83.385 ;
        RECT 117.700 73.345 117.870 83.385 ;
        RECT 119.280 73.345 119.450 83.385 ;
        RECT 130.220 83.155 130.430 86.365 ;
        RECT 130.255 82.130 130.425 83.155 ;
        RECT 130.240 81.960 130.425 82.130 ;
        RECT 125.180 80.520 125.410 81.340 ;
        RECT 124.860 80.350 126.240 80.520 ;
        RECT 126.840 80.510 127.070 81.330 ;
        RECT 126.520 80.340 127.900 80.510 ;
        RECT 127.645 79.510 127.815 79.605 ;
        RECT 126.835 79.240 127.815 79.510 ;
        RECT 127.645 78.570 127.815 79.240 ;
        RECT 126.835 78.330 127.815 78.570 ;
        RECT 127.645 78.225 127.815 78.330 ;
        RECT 127.675 77.175 127.845 78.005 ;
        RECT 126.855 76.945 127.845 77.175 ;
        RECT 127.675 76.935 127.845 76.945 ;
        RECT 127.675 76.625 127.860 76.935 ;
        RECT 125.280 75.240 125.610 75.245 ;
        RECT 125.280 75.235 127.385 75.240 ;
        RECT 127.680 75.235 127.860 76.625 ;
        RECT 125.280 75.070 127.860 75.235 ;
        RECT 125.280 75.065 125.610 75.070 ;
        RECT 125.435 75.055 125.605 75.065 ;
        RECT 127.215 75.055 127.860 75.070 ;
        RECT 127.230 75.025 127.860 75.055 ;
        RECT 127.230 75.015 127.850 75.025 ;
        RECT 22.185 53.615 33.175 53.785 ;
        RECT 22.185 46.855 22.355 53.615 ;
        RECT 33.005 46.855 33.175 53.615 ;
        RECT 35.535 53.215 35.705 53.745 ;
        RECT 36.885 53.155 37.925 53.495 ;
        RECT 104.815 53.155 105.855 53.495 ;
        RECT 107.035 53.215 107.205 53.745 ;
        RECT 109.565 53.615 120.555 53.785 ;
        RECT 35.535 49.025 35.705 49.555 ;
        RECT 36.885 49.275 37.925 49.615 ;
        RECT 104.815 49.275 105.855 49.615 ;
        RECT 107.035 49.025 107.205 49.555 ;
        RECT 22.185 46.685 33.175 46.855 ;
        RECT 37.015 46.745 37.355 47.415 ;
        RECT 105.385 46.745 105.725 47.415 ;
        RECT 109.565 46.855 109.735 53.615 ;
        RECT 120.385 46.855 120.555 53.615 ;
        RECT 109.565 46.685 120.555 46.855 ;
        RECT 23.200 42.310 23.540 42.980 ;
        RECT 27.380 42.870 38.370 43.040 ;
        RECT 22.630 40.110 23.670 40.450 ;
        RECT 24.850 40.170 25.020 40.700 ;
        RECT 15.655 39.380 15.825 39.475 ;
        RECT 15.655 39.110 16.635 39.380 ;
        RECT 15.655 38.440 15.825 39.110 ;
        RECT 15.655 38.200 16.635 38.440 ;
        RECT 15.655 38.095 15.825 38.200 ;
        RECT 12.985 37.580 13.170 37.750 ;
        RECT 12.985 37.065 13.155 37.580 ;
        RECT 14.710 37.065 15.230 37.095 ;
        RECT 12.985 36.505 15.230 37.065 ;
        RECT 12.970 36.475 15.230 36.505 ;
        RECT 12.970 36.465 15.080 36.475 ;
        RECT 12.970 33.255 13.180 36.465 ;
        RECT 22.630 36.230 23.670 36.570 ;
        RECT 24.850 35.980 25.020 36.510 ;
        RECT 27.380 36.110 27.550 42.870 ;
        RECT 28.840 36.970 29.010 42.010 ;
        RECT 30.420 36.970 30.590 42.010 ;
        RECT 32.000 36.970 32.170 42.010 ;
        RECT 33.580 36.970 33.750 42.010 ;
        RECT 35.160 36.970 35.330 42.010 ;
        RECT 36.740 36.970 36.910 42.010 ;
        RECT 38.200 36.110 38.370 42.870 ;
        RECT 27.380 35.940 38.370 36.110 ;
        RECT 104.370 42.870 115.360 43.040 ;
        RECT 104.370 36.110 104.540 42.870 ;
        RECT 105.830 36.970 106.000 42.010 ;
        RECT 107.410 36.970 107.580 42.010 ;
        RECT 108.990 36.970 109.160 42.010 ;
        RECT 110.570 36.970 110.740 42.010 ;
        RECT 112.150 36.970 112.320 42.010 ;
        RECT 113.730 36.970 113.900 42.010 ;
        RECT 115.190 36.110 115.360 42.870 ;
        RECT 119.200 42.310 119.540 42.980 ;
        RECT 117.720 40.170 117.890 40.700 ;
        RECT 119.070 40.110 120.110 40.450 ;
        RECT 126.915 39.380 127.085 39.475 ;
        RECT 126.105 39.110 127.085 39.380 ;
        RECT 126.915 38.440 127.085 39.110 ;
        RECT 126.105 38.200 127.085 38.440 ;
        RECT 126.915 38.095 127.085 38.200 ;
        RECT 129.570 37.580 129.755 37.750 ;
        RECT 127.510 37.065 128.030 37.095 ;
        RECT 129.585 37.065 129.755 37.580 ;
        RECT 104.370 35.940 115.360 36.110 ;
        RECT 117.720 35.980 117.890 36.510 ;
        RECT 119.070 36.230 120.110 36.570 ;
        RECT 127.510 36.505 129.755 37.065 ;
        RECT 127.510 36.475 129.770 36.505 ;
        RECT 127.660 36.465 129.770 36.475 ;
        RECT 16.170 34.720 16.400 35.540 ;
        RECT 17.890 34.720 18.120 35.540 ;
        RECT 124.620 34.720 124.850 35.540 ;
        RECT 126.340 34.720 126.570 35.540 ;
        RECT 15.340 34.550 16.720 34.720 ;
        RECT 17.060 34.550 18.440 34.720 ;
        RECT 124.300 34.550 125.680 34.720 ;
        RECT 126.020 34.550 127.400 34.720 ;
        RECT 12.975 32.230 13.145 33.255 ;
        RECT 12.975 32.060 13.160 32.230 ;
        RECT 16.330 30.610 16.560 31.430 ;
        RECT 17.990 30.620 18.220 31.440 ;
        RECT 15.500 30.440 16.880 30.610 ;
        RECT 17.160 30.450 18.540 30.620 ;
        RECT 15.585 29.610 15.755 29.705 ;
        RECT 15.585 29.340 16.565 29.610 ;
        RECT 15.585 28.670 15.755 29.340 ;
        RECT 15.585 28.430 16.565 28.670 ;
        RECT 15.585 28.325 15.755 28.430 ;
        RECT 15.555 27.275 15.725 28.105 ;
        RECT 15.555 27.045 16.545 27.275 ;
        RECT 15.555 27.035 15.725 27.045 ;
        RECT 15.540 26.725 15.725 27.035 ;
        RECT 15.540 25.335 15.720 26.725 ;
        RECT 17.790 25.340 18.120 25.345 ;
        RECT 16.015 25.335 18.120 25.340 ;
        RECT 15.540 25.170 18.120 25.335 ;
        RECT 15.540 25.155 16.185 25.170 ;
        RECT 17.790 25.165 18.120 25.170 ;
        RECT 17.795 25.155 17.965 25.165 ;
        RECT 15.540 25.125 16.170 25.155 ;
        RECT 15.550 25.115 16.170 25.125 ;
        RECT 23.950 23.445 24.120 33.485 ;
        RECT 25.530 23.445 25.700 33.485 ;
        RECT 27.110 23.445 27.280 33.485 ;
        RECT 28.690 23.445 28.860 33.485 ;
        RECT 30.270 23.445 30.440 33.485 ;
        RECT 31.850 23.445 32.020 33.485 ;
        RECT 33.430 23.445 33.600 33.485 ;
        RECT 35.010 23.445 35.180 33.485 ;
        RECT 36.590 23.445 36.760 33.485 ;
        RECT 105.980 23.445 106.150 33.485 ;
        RECT 107.560 23.445 107.730 33.485 ;
        RECT 109.140 23.445 109.310 33.485 ;
        RECT 110.720 23.445 110.890 33.485 ;
        RECT 112.300 23.445 112.470 33.485 ;
        RECT 113.880 23.445 114.050 33.485 ;
        RECT 115.460 23.445 115.630 33.485 ;
        RECT 117.040 23.445 117.210 33.485 ;
        RECT 118.620 23.445 118.790 33.485 ;
        RECT 129.560 33.255 129.770 36.465 ;
        RECT 129.595 32.230 129.765 33.255 ;
        RECT 129.580 32.060 129.765 32.230 ;
        RECT 124.520 30.620 124.750 31.440 ;
        RECT 124.200 30.450 125.580 30.620 ;
        RECT 126.180 30.610 126.410 31.430 ;
        RECT 125.860 30.440 127.240 30.610 ;
        RECT 126.985 29.610 127.155 29.705 ;
        RECT 126.175 29.340 127.155 29.610 ;
        RECT 126.985 28.670 127.155 29.340 ;
        RECT 126.175 28.430 127.155 28.670 ;
        RECT 126.985 28.325 127.155 28.430 ;
        RECT 127.015 27.275 127.185 28.105 ;
        RECT 126.195 27.045 127.185 27.275 ;
        RECT 127.015 27.035 127.185 27.045 ;
        RECT 127.015 26.725 127.200 27.035 ;
        RECT 124.620 25.340 124.950 25.345 ;
        RECT 124.620 25.335 126.725 25.340 ;
        RECT 127.020 25.335 127.200 26.725 ;
        RECT 124.620 25.170 127.200 25.335 ;
        RECT 124.620 25.165 124.950 25.170 ;
        RECT 124.775 25.155 124.945 25.165 ;
        RECT 126.555 25.155 127.200 25.170 ;
        RECT 126.570 25.125 127.200 25.155 ;
        RECT 126.570 25.115 127.190 25.125 ;
      LAYER met1 ;
        RECT 21.795 201.955 32.905 202.185 ;
        RECT 35.175 202.095 37.075 202.325 ;
        RECT 21.795 195.255 22.085 201.955 ;
        RECT 35.175 201.525 35.405 202.095 ;
        RECT 36.555 201.865 37.075 202.095 ;
        RECT 105.995 202.095 107.895 202.325 ;
        RECT 105.995 201.865 106.515 202.095 ;
        RECT 36.555 201.525 37.595 201.865 ;
        RECT 105.475 201.525 106.515 201.865 ;
        RECT 107.665 201.525 107.895 202.095 ;
        RECT 110.165 201.955 121.275 202.185 ;
        RECT 35.175 197.415 35.405 197.985 ;
        RECT 36.555 197.645 37.595 197.985 ;
        RECT 105.475 197.645 106.515 197.985 ;
        RECT 36.555 197.415 37.075 197.645 ;
        RECT 35.175 197.185 37.075 197.415 ;
        RECT 105.995 197.415 106.515 197.645 ;
        RECT 107.665 197.415 107.895 197.985 ;
        RECT 105.995 197.185 107.895 197.415 ;
        RECT 36.685 195.545 37.025 195.715 ;
        RECT 106.045 195.545 106.385 195.715 ;
        RECT 35.685 195.495 36.085 195.515 ;
        RECT 33.545 195.265 36.085 195.495 ;
        RECT 33.545 195.255 33.775 195.265 ;
        RECT 21.795 195.025 33.775 195.255 ;
        RECT 35.685 195.245 36.085 195.265 ;
        RECT 36.685 195.215 37.065 195.545 ;
        RECT 106.005 195.215 106.385 195.545 ;
        RECT 106.985 195.495 107.385 195.515 ;
        RECT 106.985 195.265 109.525 195.495 ;
        RECT 106.985 195.245 107.385 195.265 ;
        RECT 109.295 195.255 109.525 195.265 ;
        RECT 120.985 195.255 121.275 201.955 ;
        RECT 36.685 195.115 37.025 195.215 ;
        RECT 106.045 195.115 106.385 195.215 ;
        RECT 109.295 195.025 121.275 195.255 ;
        RECT 4.110 193.080 5.890 193.490 ;
        RECT 9.020 193.080 10.100 193.085 ;
        RECT 4.110 192.995 16.030 193.080 ;
        RECT 18.980 192.995 21.200 193.015 ;
        RECT 4.110 192.025 21.200 192.995 ;
        RECT 4.110 192.010 16.030 192.025 ;
        RECT 4.110 191.660 5.890 192.010 ;
        RECT 3.930 172.880 6.180 173.680 ;
        RECT 9.020 172.880 10.100 192.010 ;
        RECT 15.160 188.775 15.700 192.010 ;
        RECT 17.980 192.005 21.200 192.025 ;
        RECT 121.870 192.995 124.090 193.015 ;
        RECT 121.870 192.935 127.610 192.995 ;
        RECT 133.040 192.935 135.235 223.055 ;
        RECT 121.870 192.025 135.235 192.935 ;
        RECT 121.870 192.005 125.090 192.025 ;
        RECT 17.980 191.995 18.980 192.005 ;
        RECT 124.090 191.995 125.090 192.005 ;
        RECT 22.870 191.250 23.210 191.350 ;
        RECT 22.830 190.920 23.210 191.250 ;
        RECT 23.810 191.200 24.210 191.220 ;
        RECT 26.120 191.210 38.100 191.440 ;
        RECT 26.120 191.200 26.350 191.210 ;
        RECT 23.810 190.970 26.350 191.200 ;
        RECT 23.810 190.950 24.210 190.970 ;
        RECT 22.870 190.750 23.210 190.920 ;
        RECT 22.820 189.050 24.720 189.280 ;
        RECT 22.820 188.820 23.340 189.050 ;
        RECT 15.110 187.795 15.700 188.775 ;
        RECT 22.300 188.480 23.340 188.820 ;
        RECT 24.490 188.480 24.720 189.050 ;
        RECT 14.420 186.785 14.810 186.805 ;
        RECT 15.170 186.785 15.650 187.795 ;
        RECT 14.420 186.475 15.650 186.785 ;
        RECT 14.420 183.245 14.810 186.475 ;
        RECT 15.170 186.465 15.650 186.475 ;
        RECT 28.460 185.360 28.730 190.360 ;
        RECT 30.040 185.360 30.310 190.360 ;
        RECT 31.620 185.360 31.890 190.360 ;
        RECT 33.200 185.360 33.470 190.360 ;
        RECT 34.780 185.360 35.050 190.360 ;
        RECT 36.360 185.360 36.630 190.360 ;
        RECT 22.300 184.600 23.340 184.940 ;
        RECT 22.820 184.370 23.340 184.600 ;
        RECT 24.490 184.370 24.720 184.940 ;
        RECT 37.810 184.510 38.100 191.210 ;
        RECT 22.820 184.140 24.720 184.370 ;
        RECT 26.990 184.280 38.100 184.510 ;
        RECT 104.970 191.210 116.950 191.440 ;
        RECT 119.860 191.250 120.200 191.350 ;
        RECT 104.970 184.510 105.260 191.210 ;
        RECT 116.720 191.200 116.950 191.210 ;
        RECT 118.860 191.200 119.260 191.220 ;
        RECT 116.720 190.970 119.260 191.200 ;
        RECT 118.860 190.950 119.260 190.970 ;
        RECT 119.860 190.920 120.240 191.250 ;
        RECT 119.860 190.750 120.200 190.920 ;
        RECT 106.440 185.360 106.710 190.360 ;
        RECT 108.020 185.360 108.290 190.360 ;
        RECT 109.600 185.360 109.870 190.360 ;
        RECT 111.180 185.360 111.450 190.360 ;
        RECT 112.760 185.360 113.030 190.360 ;
        RECT 114.340 185.360 114.610 190.360 ;
        RECT 118.350 189.050 120.250 189.280 ;
        RECT 118.350 188.480 118.580 189.050 ;
        RECT 119.730 188.820 120.250 189.050 ;
        RECT 119.730 188.480 120.770 188.820 ;
        RECT 127.370 188.775 127.910 192.025 ;
        RECT 127.370 187.795 127.960 188.775 ;
        RECT 127.420 186.785 127.900 187.795 ;
        RECT 128.260 186.785 128.650 186.805 ;
        RECT 127.420 186.475 128.650 186.785 ;
        RECT 127.420 186.465 127.900 186.475 ;
        RECT 104.970 184.280 116.080 184.510 ;
        RECT 118.350 184.370 118.580 184.940 ;
        RECT 119.730 184.600 120.770 184.940 ;
        RECT 119.730 184.370 120.250 184.600 ;
        RECT 118.350 184.140 120.250 184.370 ;
        RECT 16.230 183.245 16.880 183.255 ;
        RECT 126.190 183.245 126.840 183.255 ;
        RECT 128.260 183.245 128.650 186.475 ;
        RECT 14.410 182.775 18.110 183.245 ;
        RECT 14.410 182.765 14.860 182.775 ;
        RECT 15.010 182.765 18.110 182.775 ;
        RECT 124.960 182.775 128.660 183.245 ;
        RECT 124.960 182.765 128.060 182.775 ;
        RECT 128.210 182.765 128.660 182.775 ;
        RECT 14.410 182.605 14.840 182.765 ;
        RECT 128.230 182.605 128.660 182.765 ;
        RECT 14.410 181.325 14.940 182.605 ;
        RECT 14.410 180.425 14.900 181.325 ;
        RECT 14.410 179.175 14.940 180.425 ;
        RECT 14.410 179.135 15.290 179.175 ;
        RECT 16.470 179.145 16.880 179.155 ;
        RECT 16.470 179.135 18.210 179.145 ;
        RECT 14.410 178.675 18.210 179.135 ;
        RECT 14.440 178.665 18.210 178.675 ;
        RECT 14.440 178.655 16.700 178.665 ;
        RECT 14.440 178.625 14.940 178.655 ;
        RECT 15.120 178.075 15.570 178.655 ;
        RECT 15.100 176.755 15.580 178.075 ;
        RECT 15.090 176.475 15.580 176.755 ;
        RECT 15.070 176.435 15.580 176.475 ;
        RECT 15.070 175.095 15.550 176.435 ;
        RECT 3.930 171.465 10.270 172.880 ;
        RECT 23.570 171.830 23.840 181.840 ;
        RECT 25.150 171.830 25.420 181.840 ;
        RECT 26.730 171.830 27.000 181.840 ;
        RECT 28.310 171.830 28.580 181.840 ;
        RECT 29.890 171.830 30.160 181.840 ;
        RECT 31.470 171.830 31.740 181.840 ;
        RECT 33.050 171.830 33.320 181.840 ;
        RECT 34.630 171.830 34.900 181.840 ;
        RECT 36.210 171.830 36.480 181.840 ;
        RECT 106.590 171.830 106.860 181.840 ;
        RECT 108.170 171.830 108.440 181.840 ;
        RECT 109.750 171.830 110.020 181.840 ;
        RECT 111.330 171.830 111.600 181.840 ;
        RECT 112.910 171.830 113.180 181.840 ;
        RECT 114.490 171.830 114.760 181.840 ;
        RECT 116.070 171.830 116.340 181.840 ;
        RECT 117.650 171.830 117.920 181.840 ;
        RECT 119.230 171.830 119.500 181.840 ;
        RECT 128.130 181.325 128.660 182.605 ;
        RECT 128.170 180.425 128.660 181.325 ;
        RECT 128.130 179.175 128.660 180.425 ;
        RECT 126.190 179.145 126.600 179.155 ;
        RECT 124.860 179.135 126.600 179.145 ;
        RECT 127.780 179.135 128.660 179.175 ;
        RECT 124.860 178.675 128.660 179.135 ;
        RECT 124.860 178.665 128.630 178.675 ;
        RECT 126.370 178.655 128.630 178.665 ;
        RECT 127.500 178.075 127.950 178.655 ;
        RECT 128.130 178.625 128.630 178.655 ;
        RECT 127.490 176.755 127.970 178.075 ;
        RECT 127.490 176.475 127.980 176.755 ;
        RECT 127.490 176.435 128.000 176.475 ;
        RECT 127.520 175.095 128.000 176.435 ;
        RECT 3.930 170.970 6.180 171.465 ;
        RECT 9.020 143.340 10.100 171.465 ;
        RECT 21.795 152.385 32.905 152.615 ;
        RECT 35.175 152.525 37.075 152.755 ;
        RECT 21.795 145.685 22.085 152.385 ;
        RECT 35.175 151.955 35.405 152.525 ;
        RECT 36.555 152.295 37.075 152.525 ;
        RECT 105.995 152.525 107.895 152.755 ;
        RECT 105.995 152.295 106.515 152.525 ;
        RECT 36.555 151.955 37.595 152.295 ;
        RECT 105.475 151.955 106.515 152.295 ;
        RECT 107.665 151.955 107.895 152.525 ;
        RECT 110.165 152.385 121.275 152.615 ;
        RECT 35.175 147.845 35.405 148.415 ;
        RECT 36.555 148.075 37.595 148.415 ;
        RECT 105.475 148.075 106.515 148.415 ;
        RECT 36.555 147.845 37.075 148.075 ;
        RECT 35.175 147.615 37.075 147.845 ;
        RECT 105.995 147.845 106.515 148.075 ;
        RECT 107.665 147.845 107.895 148.415 ;
        RECT 105.995 147.615 107.895 147.845 ;
        RECT 36.685 145.975 37.025 146.145 ;
        RECT 106.045 145.975 106.385 146.145 ;
        RECT 35.685 145.925 36.085 145.945 ;
        RECT 33.545 145.695 36.085 145.925 ;
        RECT 33.545 145.685 33.775 145.695 ;
        RECT 21.795 145.455 33.775 145.685 ;
        RECT 35.685 145.675 36.085 145.695 ;
        RECT 36.685 145.645 37.065 145.975 ;
        RECT 106.005 145.645 106.385 145.975 ;
        RECT 106.985 145.925 107.385 145.945 ;
        RECT 106.985 145.695 109.525 145.925 ;
        RECT 106.985 145.675 107.385 145.695 ;
        RECT 109.295 145.685 109.525 145.695 ;
        RECT 120.985 145.685 121.275 152.385 ;
        RECT 36.685 145.545 37.025 145.645 ;
        RECT 106.045 145.545 106.385 145.645 ;
        RECT 109.295 145.455 121.275 145.685 ;
        RECT 18.980 143.425 21.200 143.445 ;
        RECT 15.460 143.365 21.200 143.425 ;
        RECT 15.160 143.340 21.200 143.365 ;
        RECT 9.020 142.455 21.200 143.340 ;
        RECT 9.020 142.260 16.590 142.455 ;
        RECT 17.980 142.435 21.200 142.455 ;
        RECT 121.870 143.425 124.090 143.445 ;
        RECT 133.040 143.425 135.235 192.025 ;
        RECT 121.870 142.455 135.235 143.425 ;
        RECT 121.870 142.435 125.090 142.455 ;
        RECT 17.980 142.425 18.980 142.435 ;
        RECT 124.090 142.425 125.090 142.435 ;
        RECT 9.030 115.400 10.090 142.260 ;
        RECT 15.160 139.205 15.700 142.260 ;
        RECT 22.870 141.680 23.210 141.780 ;
        RECT 22.830 141.350 23.210 141.680 ;
        RECT 23.810 141.630 24.210 141.650 ;
        RECT 26.120 141.640 38.100 141.870 ;
        RECT 26.120 141.630 26.350 141.640 ;
        RECT 23.810 141.400 26.350 141.630 ;
        RECT 23.810 141.380 24.210 141.400 ;
        RECT 22.870 141.180 23.210 141.350 ;
        RECT 22.820 139.480 24.720 139.710 ;
        RECT 22.820 139.250 23.340 139.480 ;
        RECT 15.110 138.225 15.700 139.205 ;
        RECT 22.300 138.910 23.340 139.250 ;
        RECT 24.490 138.910 24.720 139.480 ;
        RECT 14.420 137.215 14.810 137.235 ;
        RECT 15.170 137.215 15.650 138.225 ;
        RECT 14.420 136.905 15.650 137.215 ;
        RECT 14.420 133.675 14.810 136.905 ;
        RECT 15.170 136.895 15.650 136.905 ;
        RECT 28.460 135.790 28.730 140.790 ;
        RECT 30.040 135.790 30.310 140.790 ;
        RECT 31.620 135.790 31.890 140.790 ;
        RECT 33.200 135.790 33.470 140.790 ;
        RECT 34.780 135.790 35.050 140.790 ;
        RECT 36.360 135.790 36.630 140.790 ;
        RECT 22.300 135.030 23.340 135.370 ;
        RECT 22.820 134.800 23.340 135.030 ;
        RECT 24.490 134.800 24.720 135.370 ;
        RECT 37.810 134.940 38.100 141.640 ;
        RECT 22.820 134.570 24.720 134.800 ;
        RECT 26.990 134.710 38.100 134.940 ;
        RECT 104.970 141.640 116.950 141.870 ;
        RECT 119.860 141.680 120.200 141.780 ;
        RECT 104.970 134.940 105.260 141.640 ;
        RECT 116.720 141.630 116.950 141.640 ;
        RECT 118.860 141.630 119.260 141.650 ;
        RECT 116.720 141.400 119.260 141.630 ;
        RECT 118.860 141.380 119.260 141.400 ;
        RECT 119.860 141.350 120.240 141.680 ;
        RECT 119.860 141.180 120.200 141.350 ;
        RECT 106.440 135.790 106.710 140.790 ;
        RECT 108.020 135.790 108.290 140.790 ;
        RECT 109.600 135.790 109.870 140.790 ;
        RECT 111.180 135.790 111.450 140.790 ;
        RECT 112.760 135.790 113.030 140.790 ;
        RECT 114.340 135.790 114.610 140.790 ;
        RECT 118.350 139.480 120.250 139.710 ;
        RECT 118.350 138.910 118.580 139.480 ;
        RECT 119.730 139.250 120.250 139.480 ;
        RECT 119.730 138.910 120.770 139.250 ;
        RECT 127.370 139.205 127.910 142.455 ;
        RECT 127.370 138.225 127.960 139.205 ;
        RECT 127.420 137.215 127.900 138.225 ;
        RECT 128.260 137.215 128.650 137.235 ;
        RECT 127.420 136.905 128.650 137.215 ;
        RECT 127.420 136.895 127.900 136.905 ;
        RECT 104.970 134.710 116.080 134.940 ;
        RECT 118.350 134.800 118.580 135.370 ;
        RECT 119.730 135.030 120.770 135.370 ;
        RECT 119.730 134.800 120.250 135.030 ;
        RECT 118.350 134.570 120.250 134.800 ;
        RECT 16.230 133.675 16.880 133.685 ;
        RECT 126.190 133.675 126.840 133.685 ;
        RECT 128.260 133.675 128.650 136.905 ;
        RECT 14.410 133.205 18.110 133.675 ;
        RECT 14.410 133.195 14.860 133.205 ;
        RECT 15.010 133.195 18.110 133.205 ;
        RECT 124.960 133.205 128.660 133.675 ;
        RECT 124.960 133.195 128.060 133.205 ;
        RECT 128.210 133.195 128.660 133.205 ;
        RECT 14.410 133.035 14.840 133.195 ;
        RECT 128.230 133.035 128.660 133.195 ;
        RECT 14.410 131.755 14.940 133.035 ;
        RECT 14.410 130.855 14.900 131.755 ;
        RECT 14.410 129.605 14.940 130.855 ;
        RECT 14.410 129.565 15.290 129.605 ;
        RECT 16.470 129.575 16.880 129.585 ;
        RECT 16.470 129.565 18.210 129.575 ;
        RECT 14.410 129.105 18.210 129.565 ;
        RECT 14.440 129.095 18.210 129.105 ;
        RECT 14.440 129.085 16.700 129.095 ;
        RECT 14.440 129.055 14.940 129.085 ;
        RECT 15.120 128.505 15.570 129.085 ;
        RECT 15.100 127.185 15.580 128.505 ;
        RECT 15.090 126.905 15.580 127.185 ;
        RECT 15.070 126.865 15.580 126.905 ;
        RECT 15.070 125.525 15.550 126.865 ;
        RECT 23.570 122.260 23.840 132.270 ;
        RECT 25.150 122.260 25.420 132.270 ;
        RECT 26.730 122.260 27.000 132.270 ;
        RECT 28.310 122.260 28.580 132.270 ;
        RECT 29.890 122.260 30.160 132.270 ;
        RECT 31.470 122.260 31.740 132.270 ;
        RECT 33.050 122.260 33.320 132.270 ;
        RECT 34.630 122.260 34.900 132.270 ;
        RECT 36.210 122.260 36.480 132.270 ;
        RECT 106.590 122.260 106.860 132.270 ;
        RECT 108.170 122.260 108.440 132.270 ;
        RECT 109.750 122.260 110.020 132.270 ;
        RECT 111.330 122.260 111.600 132.270 ;
        RECT 112.910 122.260 113.180 132.270 ;
        RECT 114.490 122.260 114.760 132.270 ;
        RECT 116.070 122.260 116.340 132.270 ;
        RECT 117.650 122.260 117.920 132.270 ;
        RECT 119.230 122.260 119.500 132.270 ;
        RECT 128.130 131.755 128.660 133.035 ;
        RECT 128.170 130.855 128.660 131.755 ;
        RECT 128.130 129.605 128.660 130.855 ;
        RECT 126.190 129.575 126.600 129.585 ;
        RECT 124.860 129.565 126.600 129.575 ;
        RECT 127.780 129.565 128.660 129.605 ;
        RECT 124.860 129.105 128.660 129.565 ;
        RECT 124.860 129.095 128.630 129.105 ;
        RECT 126.370 129.085 128.630 129.095 ;
        RECT 127.500 128.505 127.950 129.085 ;
        RECT 128.130 129.055 128.630 129.085 ;
        RECT 127.490 127.185 127.970 128.505 ;
        RECT 127.490 126.905 127.980 127.185 ;
        RECT 127.490 126.865 128.000 126.905 ;
        RECT 127.520 125.525 128.000 126.865 ;
        RECT 3.990 114.530 6.210 115.330 ;
        RECT 9.030 114.530 10.130 115.400 ;
        RECT 3.990 113.115 10.250 114.530 ;
        RECT 3.990 112.620 6.210 113.115 ;
        RECT 9.030 112.600 10.130 113.115 ;
        RECT 9.030 103.450 10.090 112.600 ;
        RECT 22.455 104.155 33.565 104.385 ;
        RECT 35.835 104.295 37.735 104.525 ;
        RECT 9.030 101.970 10.150 103.450 ;
        RECT 9.030 95.180 10.090 101.970 ;
        RECT 22.455 97.455 22.745 104.155 ;
        RECT 35.835 103.725 36.065 104.295 ;
        RECT 37.215 104.065 37.735 104.295 ;
        RECT 37.215 103.725 38.255 104.065 ;
        RECT 105.995 103.625 107.895 103.855 ;
        RECT 105.995 103.395 106.515 103.625 ;
        RECT 105.475 103.055 106.515 103.395 ;
        RECT 107.665 103.055 107.895 103.625 ;
        RECT 110.165 103.485 121.275 103.715 ;
        RECT 35.835 99.615 36.065 100.185 ;
        RECT 37.215 99.845 38.255 100.185 ;
        RECT 37.215 99.615 37.735 99.845 ;
        RECT 35.835 99.385 37.735 99.615 ;
        RECT 105.475 99.175 106.515 99.515 ;
        RECT 105.995 98.945 106.515 99.175 ;
        RECT 107.665 98.945 107.895 99.515 ;
        RECT 105.995 98.715 107.895 98.945 ;
        RECT 37.345 97.745 37.685 97.915 ;
        RECT 36.345 97.695 36.745 97.715 ;
        RECT 34.205 97.465 36.745 97.695 ;
        RECT 34.205 97.455 34.435 97.465 ;
        RECT 22.455 97.225 34.435 97.455 ;
        RECT 36.345 97.445 36.745 97.465 ;
        RECT 37.345 97.415 37.725 97.745 ;
        RECT 37.345 97.315 37.685 97.415 ;
        RECT 106.045 97.075 106.385 97.245 ;
        RECT 106.005 96.745 106.385 97.075 ;
        RECT 106.985 97.025 107.385 97.045 ;
        RECT 106.985 96.795 109.525 97.025 ;
        RECT 106.985 96.775 107.385 96.795 ;
        RECT 109.295 96.785 109.525 96.795 ;
        RECT 120.985 96.785 121.275 103.485 ;
        RECT 106.045 96.645 106.385 96.745 ;
        RECT 109.295 96.555 121.275 96.785 ;
        RECT 19.640 95.195 21.860 95.215 ;
        RECT 16.120 95.180 21.860 95.195 ;
        RECT 9.030 94.225 21.860 95.180 ;
        RECT 9.030 94.120 17.110 94.225 ;
        RECT 18.640 94.205 21.860 94.225 ;
        RECT 121.870 94.525 124.090 94.545 ;
        RECT 133.040 94.525 135.235 142.455 ;
        RECT 18.640 94.195 19.640 94.205 ;
        RECT 9.045 69.170 10.080 94.120 ;
        RECT 15.820 90.975 16.360 94.120 ;
        RECT 23.530 93.450 23.870 93.550 ;
        RECT 23.490 93.120 23.870 93.450 ;
        RECT 24.470 93.400 24.870 93.420 ;
        RECT 26.780 93.410 38.760 93.640 ;
        RECT 121.870 93.555 135.235 94.525 ;
        RECT 121.870 93.535 125.090 93.555 ;
        RECT 124.090 93.525 125.090 93.535 ;
        RECT 26.780 93.400 27.010 93.410 ;
        RECT 24.470 93.170 27.010 93.400 ;
        RECT 24.470 93.150 24.870 93.170 ;
        RECT 23.530 92.950 23.870 93.120 ;
        RECT 23.480 91.250 25.380 91.480 ;
        RECT 23.480 91.020 24.000 91.250 ;
        RECT 15.770 89.995 16.360 90.975 ;
        RECT 22.960 90.680 24.000 91.020 ;
        RECT 25.150 90.680 25.380 91.250 ;
        RECT 15.080 88.985 15.470 89.005 ;
        RECT 15.830 88.985 16.310 89.995 ;
        RECT 15.080 88.675 16.310 88.985 ;
        RECT 15.080 85.445 15.470 88.675 ;
        RECT 15.830 88.665 16.310 88.675 ;
        RECT 29.120 87.560 29.390 92.560 ;
        RECT 30.700 87.560 30.970 92.560 ;
        RECT 32.280 87.560 32.550 92.560 ;
        RECT 33.860 87.560 34.130 92.560 ;
        RECT 35.440 87.560 35.710 92.560 ;
        RECT 37.020 87.560 37.290 92.560 ;
        RECT 22.960 86.800 24.000 87.140 ;
        RECT 23.480 86.570 24.000 86.800 ;
        RECT 25.150 86.570 25.380 87.140 ;
        RECT 38.470 86.710 38.760 93.410 ;
        RECT 23.480 86.340 25.380 86.570 ;
        RECT 27.650 86.480 38.760 86.710 ;
        RECT 104.970 92.740 116.950 92.970 ;
        RECT 119.860 92.780 120.200 92.880 ;
        RECT 104.970 86.040 105.260 92.740 ;
        RECT 116.720 92.730 116.950 92.740 ;
        RECT 118.860 92.730 119.260 92.750 ;
        RECT 116.720 92.500 119.260 92.730 ;
        RECT 118.860 92.480 119.260 92.500 ;
        RECT 119.860 92.450 120.240 92.780 ;
        RECT 119.860 92.280 120.200 92.450 ;
        RECT 106.440 86.890 106.710 91.890 ;
        RECT 108.020 86.890 108.290 91.890 ;
        RECT 109.600 86.890 109.870 91.890 ;
        RECT 111.180 86.890 111.450 91.890 ;
        RECT 112.760 86.890 113.030 91.890 ;
        RECT 114.340 86.890 114.610 91.890 ;
        RECT 118.350 90.580 120.250 90.810 ;
        RECT 118.350 90.010 118.580 90.580 ;
        RECT 119.730 90.350 120.250 90.580 ;
        RECT 119.730 90.010 120.770 90.350 ;
        RECT 127.370 90.305 127.910 93.555 ;
        RECT 127.370 89.325 127.960 90.305 ;
        RECT 127.420 88.315 127.900 89.325 ;
        RECT 128.260 88.315 128.650 88.335 ;
        RECT 127.420 88.005 128.650 88.315 ;
        RECT 127.420 87.995 127.900 88.005 ;
        RECT 104.970 85.810 116.080 86.040 ;
        RECT 118.350 85.900 118.580 86.470 ;
        RECT 119.730 86.130 120.770 86.470 ;
        RECT 119.730 85.900 120.250 86.130 ;
        RECT 118.350 85.670 120.250 85.900 ;
        RECT 16.890 85.445 17.540 85.455 ;
        RECT 15.070 84.975 18.770 85.445 ;
        RECT 15.070 84.965 15.520 84.975 ;
        RECT 15.670 84.965 18.770 84.975 ;
        RECT 15.070 84.805 15.500 84.965 ;
        RECT 15.070 83.525 15.600 84.805 ;
        RECT 126.190 84.775 126.840 84.785 ;
        RECT 128.260 84.775 128.650 88.005 ;
        RECT 124.960 84.305 128.660 84.775 ;
        RECT 124.960 84.295 128.060 84.305 ;
        RECT 128.210 84.295 128.660 84.305 ;
        RECT 128.230 84.135 128.660 84.295 ;
        RECT 15.070 82.625 15.560 83.525 ;
        RECT 15.070 81.375 15.600 82.625 ;
        RECT 15.070 81.335 15.950 81.375 ;
        RECT 17.130 81.345 17.540 81.355 ;
        RECT 17.130 81.335 18.870 81.345 ;
        RECT 15.070 80.875 18.870 81.335 ;
        RECT 15.100 80.865 18.870 80.875 ;
        RECT 15.100 80.855 17.360 80.865 ;
        RECT 15.100 80.825 15.600 80.855 ;
        RECT 15.780 80.275 16.230 80.855 ;
        RECT 15.760 78.955 16.240 80.275 ;
        RECT 15.750 78.675 16.240 78.955 ;
        RECT 15.730 78.635 16.240 78.675 ;
        RECT 15.730 77.295 16.210 78.635 ;
        RECT 24.230 74.030 24.500 84.040 ;
        RECT 25.810 74.030 26.080 84.040 ;
        RECT 27.390 74.030 27.660 84.040 ;
        RECT 28.970 74.030 29.240 84.040 ;
        RECT 30.550 74.030 30.820 84.040 ;
        RECT 32.130 74.030 32.400 84.040 ;
        RECT 33.710 74.030 33.980 84.040 ;
        RECT 35.290 74.030 35.560 84.040 ;
        RECT 36.870 74.030 37.140 84.040 ;
        RECT 106.590 73.360 106.860 83.370 ;
        RECT 108.170 73.360 108.440 83.370 ;
        RECT 109.750 73.360 110.020 83.370 ;
        RECT 111.330 73.360 111.600 83.370 ;
        RECT 112.910 73.360 113.180 83.370 ;
        RECT 114.490 73.360 114.760 83.370 ;
        RECT 116.070 73.360 116.340 83.370 ;
        RECT 117.650 73.360 117.920 83.370 ;
        RECT 119.230 73.360 119.500 83.370 ;
        RECT 128.130 82.855 128.660 84.135 ;
        RECT 128.170 81.955 128.660 82.855 ;
        RECT 128.130 80.705 128.660 81.955 ;
        RECT 126.190 80.675 126.600 80.685 ;
        RECT 124.860 80.665 126.600 80.675 ;
        RECT 127.780 80.665 128.660 80.705 ;
        RECT 124.860 80.205 128.660 80.665 ;
        RECT 124.860 80.195 128.630 80.205 ;
        RECT 126.370 80.185 128.630 80.195 ;
        RECT 127.500 79.605 127.950 80.185 ;
        RECT 128.130 80.155 128.630 80.185 ;
        RECT 127.490 78.285 127.970 79.605 ;
        RECT 127.490 78.005 127.980 78.285 ;
        RECT 127.490 77.965 128.000 78.005 ;
        RECT 127.520 76.625 128.000 77.965 ;
        RECT 9.030 67.690 10.110 69.170 ;
        RECT 9.045 63.370 10.080 67.690 ;
        RECT 3.960 62.500 6.180 63.300 ;
        RECT 9.020 62.500 10.100 63.370 ;
        RECT 3.960 61.085 10.220 62.500 ;
        RECT 3.960 60.590 6.180 61.085 ;
        RECT 9.020 60.570 10.100 61.085 ;
        RECT 9.045 44.855 10.080 60.570 ;
        RECT 22.125 53.585 33.235 53.815 ;
        RECT 35.505 53.725 37.405 53.955 ;
        RECT 22.125 46.885 22.415 53.585 ;
        RECT 35.505 53.155 35.735 53.725 ;
        RECT 36.885 53.495 37.405 53.725 ;
        RECT 105.335 53.725 107.235 53.955 ;
        RECT 105.335 53.495 105.855 53.725 ;
        RECT 36.885 53.155 37.925 53.495 ;
        RECT 104.815 53.155 105.855 53.495 ;
        RECT 107.005 53.155 107.235 53.725 ;
        RECT 109.505 53.585 120.615 53.815 ;
        RECT 35.505 49.045 35.735 49.615 ;
        RECT 36.885 49.275 37.925 49.615 ;
        RECT 104.815 49.275 105.855 49.615 ;
        RECT 36.885 49.045 37.405 49.275 ;
        RECT 35.505 48.815 37.405 49.045 ;
        RECT 105.335 49.045 105.855 49.275 ;
        RECT 107.005 49.045 107.235 49.615 ;
        RECT 105.335 48.815 107.235 49.045 ;
        RECT 37.015 47.175 37.355 47.345 ;
        RECT 105.385 47.175 105.725 47.345 ;
        RECT 36.015 47.125 36.415 47.145 ;
        RECT 33.875 46.895 36.415 47.125 ;
        RECT 33.875 46.885 34.105 46.895 ;
        RECT 22.125 46.655 34.105 46.885 ;
        RECT 36.015 46.875 36.415 46.895 ;
        RECT 37.015 46.845 37.395 47.175 ;
        RECT 105.345 46.845 105.725 47.175 ;
        RECT 106.325 47.125 106.725 47.145 ;
        RECT 106.325 46.895 108.865 47.125 ;
        RECT 106.325 46.875 106.725 46.895 ;
        RECT 108.635 46.885 108.865 46.895 ;
        RECT 120.325 46.885 120.615 53.585 ;
        RECT 37.015 46.745 37.355 46.845 ;
        RECT 105.385 46.745 105.725 46.845 ;
        RECT 108.635 46.655 120.615 46.885 ;
        RECT 8.830 44.610 10.290 44.855 ;
        RECT 19.310 44.625 21.530 44.645 ;
        RECT 15.790 44.610 21.530 44.625 ;
        RECT 8.830 43.655 21.530 44.610 ;
        RECT 8.830 43.575 16.865 43.655 ;
        RECT 18.310 43.635 21.530 43.655 ;
        RECT 121.210 44.625 123.430 44.645 ;
        RECT 133.040 44.625 135.235 93.555 ;
        RECT 121.210 43.655 135.235 44.625 ;
        RECT 121.210 43.635 124.430 43.655 ;
        RECT 18.310 43.625 19.310 43.635 ;
        RECT 123.430 43.625 124.430 43.635 ;
        RECT 8.830 13.355 10.290 43.575 ;
        RECT 15.490 40.405 16.030 43.575 ;
        RECT 23.200 42.880 23.540 42.980 ;
        RECT 23.160 42.550 23.540 42.880 ;
        RECT 24.140 42.830 24.540 42.850 ;
        RECT 26.450 42.840 38.430 43.070 ;
        RECT 26.450 42.830 26.680 42.840 ;
        RECT 24.140 42.600 26.680 42.830 ;
        RECT 24.140 42.580 24.540 42.600 ;
        RECT 23.200 42.380 23.540 42.550 ;
        RECT 23.150 40.680 25.050 40.910 ;
        RECT 23.150 40.450 23.670 40.680 ;
        RECT 15.440 39.425 16.030 40.405 ;
        RECT 22.630 40.110 23.670 40.450 ;
        RECT 24.820 40.110 25.050 40.680 ;
        RECT 14.750 38.415 15.140 38.435 ;
        RECT 15.500 38.415 15.980 39.425 ;
        RECT 14.750 38.105 15.980 38.415 ;
        RECT 14.750 34.875 15.140 38.105 ;
        RECT 15.500 38.095 15.980 38.105 ;
        RECT 28.790 36.990 29.060 41.990 ;
        RECT 30.370 36.990 30.640 41.990 ;
        RECT 31.950 36.990 32.220 41.990 ;
        RECT 33.530 36.990 33.800 41.990 ;
        RECT 35.110 36.990 35.380 41.990 ;
        RECT 36.690 36.990 36.960 41.990 ;
        RECT 22.630 36.230 23.670 36.570 ;
        RECT 23.150 36.000 23.670 36.230 ;
        RECT 24.820 36.000 25.050 36.570 ;
        RECT 38.140 36.140 38.430 42.840 ;
        RECT 23.150 35.770 25.050 36.000 ;
        RECT 27.320 35.910 38.430 36.140 ;
        RECT 104.310 42.840 116.290 43.070 ;
        RECT 119.200 42.880 119.540 42.980 ;
        RECT 104.310 36.140 104.600 42.840 ;
        RECT 116.060 42.830 116.290 42.840 ;
        RECT 118.200 42.830 118.600 42.850 ;
        RECT 116.060 42.600 118.600 42.830 ;
        RECT 118.200 42.580 118.600 42.600 ;
        RECT 119.200 42.550 119.580 42.880 ;
        RECT 119.200 42.380 119.540 42.550 ;
        RECT 105.780 36.990 106.050 41.990 ;
        RECT 107.360 36.990 107.630 41.990 ;
        RECT 108.940 36.990 109.210 41.990 ;
        RECT 110.520 36.990 110.790 41.990 ;
        RECT 112.100 36.990 112.370 41.990 ;
        RECT 113.680 36.990 113.950 41.990 ;
        RECT 117.690 40.680 119.590 40.910 ;
        RECT 117.690 40.110 117.920 40.680 ;
        RECT 119.070 40.450 119.590 40.680 ;
        RECT 119.070 40.110 120.110 40.450 ;
        RECT 126.710 40.405 127.250 43.655 ;
        RECT 126.710 39.425 127.300 40.405 ;
        RECT 126.760 38.415 127.240 39.425 ;
        RECT 127.600 38.415 127.990 38.435 ;
        RECT 126.760 38.105 127.990 38.415 ;
        RECT 126.760 38.095 127.240 38.105 ;
        RECT 104.310 35.910 115.420 36.140 ;
        RECT 117.690 36.000 117.920 36.570 ;
        RECT 119.070 36.230 120.110 36.570 ;
        RECT 119.070 36.000 119.590 36.230 ;
        RECT 117.690 35.770 119.590 36.000 ;
        RECT 16.560 34.875 17.210 34.885 ;
        RECT 125.530 34.875 126.180 34.885 ;
        RECT 127.600 34.875 127.990 38.105 ;
        RECT 14.740 34.405 18.440 34.875 ;
        RECT 14.740 34.395 15.190 34.405 ;
        RECT 15.340 34.395 18.440 34.405 ;
        RECT 124.300 34.405 128.000 34.875 ;
        RECT 124.300 34.395 127.400 34.405 ;
        RECT 127.550 34.395 128.000 34.405 ;
        RECT 14.740 34.235 15.170 34.395 ;
        RECT 127.570 34.235 128.000 34.395 ;
        RECT 14.740 32.955 15.270 34.235 ;
        RECT 14.740 32.055 15.230 32.955 ;
        RECT 14.740 30.805 15.270 32.055 ;
        RECT 14.740 30.765 15.620 30.805 ;
        RECT 16.800 30.775 17.210 30.785 ;
        RECT 16.800 30.765 18.540 30.775 ;
        RECT 14.740 30.305 18.540 30.765 ;
        RECT 14.770 30.295 18.540 30.305 ;
        RECT 14.770 30.285 17.030 30.295 ;
        RECT 14.770 30.255 15.270 30.285 ;
        RECT 15.450 29.705 15.900 30.285 ;
        RECT 15.430 28.385 15.910 29.705 ;
        RECT 15.420 28.105 15.910 28.385 ;
        RECT 15.400 28.065 15.910 28.105 ;
        RECT 15.400 26.725 15.880 28.065 ;
        RECT 23.900 23.460 24.170 33.470 ;
        RECT 25.480 23.460 25.750 33.470 ;
        RECT 27.060 23.460 27.330 33.470 ;
        RECT 28.640 23.460 28.910 33.470 ;
        RECT 30.220 23.460 30.490 33.470 ;
        RECT 31.800 23.460 32.070 33.470 ;
        RECT 33.380 23.460 33.650 33.470 ;
        RECT 34.960 23.460 35.230 33.470 ;
        RECT 36.540 23.460 36.810 33.470 ;
        RECT 105.930 23.460 106.200 33.470 ;
        RECT 107.510 23.460 107.780 33.470 ;
        RECT 109.090 23.460 109.360 33.470 ;
        RECT 110.670 23.460 110.940 33.470 ;
        RECT 112.250 23.460 112.520 33.470 ;
        RECT 113.830 23.460 114.100 33.470 ;
        RECT 115.410 23.460 115.680 33.470 ;
        RECT 116.990 23.460 117.260 33.470 ;
        RECT 118.570 23.460 118.840 33.470 ;
        RECT 127.470 32.955 128.000 34.235 ;
        RECT 127.510 32.055 128.000 32.955 ;
        RECT 127.470 30.805 128.000 32.055 ;
        RECT 125.530 30.775 125.940 30.785 ;
        RECT 124.200 30.765 125.940 30.775 ;
        RECT 127.120 30.765 128.000 30.805 ;
        RECT 124.200 30.305 128.000 30.765 ;
        RECT 124.200 30.295 127.970 30.305 ;
        RECT 125.710 30.285 127.970 30.295 ;
        RECT 126.840 29.705 127.290 30.285 ;
        RECT 127.470 30.255 127.970 30.285 ;
        RECT 126.830 28.385 127.310 29.705 ;
        RECT 126.830 28.105 127.320 28.385 ;
        RECT 126.830 28.065 127.340 28.105 ;
        RECT 126.860 26.725 127.340 28.065 ;
        RECT 133.040 13.355 135.235 43.655 ;
        RECT 8.490 11.210 135.235 13.355 ;
        RECT 133.040 11.185 135.235 11.210 ;
      LAYER met2 ;
        RECT 36.555 201.525 37.075 202.325 ;
        RECT 105.995 201.525 106.515 202.325 ;
        RECT 36.555 197.185 37.075 197.985 ;
        RECT 105.995 197.185 106.515 197.985 ;
        RECT 35.695 195.215 36.075 195.545 ;
        RECT 36.705 195.215 37.085 195.545 ;
        RECT 105.985 195.215 106.365 195.545 ;
        RECT 106.995 195.215 107.375 195.545 ;
        RECT 4.160 191.770 5.670 193.190 ;
        RECT 20.240 192.865 20.870 192.895 ;
        RECT 20.220 192.165 20.870 192.865 ;
        RECT 122.200 192.865 122.830 192.895 ;
        RECT 122.200 192.165 122.850 192.865 ;
        RECT 20.220 192.135 20.850 192.165 ;
        RECT 122.220 192.135 122.850 192.165 ;
        RECT 22.810 190.920 23.190 191.250 ;
        RECT 23.820 190.920 24.200 191.250 ;
        RECT 118.870 190.920 119.250 191.250 ;
        RECT 119.880 190.920 120.260 191.250 ;
        RECT 22.820 188.480 23.340 189.280 ;
        RECT 119.730 188.480 120.250 189.280 ;
        RECT 28.460 185.360 36.630 187.360 ;
        RECT 106.440 185.360 114.610 187.360 ;
        RECT 22.820 184.140 23.340 184.940 ;
        RECT 119.730 184.140 120.250 184.940 ;
        RECT 20.820 179.840 36.480 181.840 ;
        RECT 106.590 179.840 122.250 181.840 ;
        RECT 20.820 176.500 22.280 179.840 ;
        RECT 120.790 176.500 122.250 179.840 ;
        RECT 20.820 174.500 36.480 176.500 ;
        RECT 106.590 174.500 122.250 176.500 ;
        RECT 4.130 171.350 5.780 173.140 ;
        RECT 36.555 151.955 37.075 152.755 ;
        RECT 105.995 151.955 106.515 152.755 ;
        RECT 36.555 147.615 37.075 148.415 ;
        RECT 105.995 147.615 106.515 148.415 ;
        RECT 35.695 145.645 36.075 145.975 ;
        RECT 36.705 145.645 37.085 145.975 ;
        RECT 105.985 145.645 106.365 145.975 ;
        RECT 106.995 145.645 107.375 145.975 ;
        RECT 20.240 143.295 20.870 143.325 ;
        RECT 20.220 142.595 20.870 143.295 ;
        RECT 122.200 143.295 122.830 143.325 ;
        RECT 122.200 142.595 122.850 143.295 ;
        RECT 20.220 142.565 20.850 142.595 ;
        RECT 122.220 142.565 122.850 142.595 ;
        RECT 22.810 141.350 23.190 141.680 ;
        RECT 23.820 141.350 24.200 141.680 ;
        RECT 118.870 141.350 119.250 141.680 ;
        RECT 119.880 141.350 120.260 141.680 ;
        RECT 22.820 138.910 23.340 139.710 ;
        RECT 119.730 138.910 120.250 139.710 ;
        RECT 28.460 135.790 36.630 137.790 ;
        RECT 106.440 135.790 114.610 137.790 ;
        RECT 22.820 134.570 23.340 135.370 ;
        RECT 119.730 134.570 120.250 135.370 ;
        RECT 20.820 130.270 36.480 132.270 ;
        RECT 106.590 130.270 122.250 132.270 ;
        RECT 20.820 126.930 22.280 130.270 ;
        RECT 120.790 126.930 122.250 130.270 ;
        RECT 20.820 124.930 36.480 126.930 ;
        RECT 106.590 124.930 122.250 126.930 ;
        RECT 4.160 113.000 5.810 114.790 ;
        RECT 37.215 103.725 37.735 104.525 ;
        RECT 105.995 103.055 106.515 103.855 ;
        RECT 37.215 99.385 37.735 100.185 ;
        RECT 105.995 98.715 106.515 99.515 ;
        RECT 36.355 97.415 36.735 97.745 ;
        RECT 37.365 97.415 37.745 97.745 ;
        RECT 105.985 96.745 106.365 97.075 ;
        RECT 106.995 96.745 107.375 97.075 ;
        RECT 20.900 95.065 21.530 95.095 ;
        RECT 20.880 94.365 21.530 95.065 ;
        RECT 122.200 94.395 122.830 94.425 ;
        RECT 20.880 94.335 21.510 94.365 ;
        RECT 122.200 93.695 122.850 94.395 ;
        RECT 122.220 93.665 122.850 93.695 ;
        RECT 23.470 93.120 23.850 93.450 ;
        RECT 24.480 93.120 24.860 93.450 ;
        RECT 118.870 92.450 119.250 92.780 ;
        RECT 119.880 92.450 120.260 92.780 ;
        RECT 23.480 90.680 24.000 91.480 ;
        RECT 119.730 90.010 120.250 90.810 ;
        RECT 29.120 87.560 37.290 89.560 ;
        RECT 23.480 86.340 24.000 87.140 ;
        RECT 106.440 86.890 114.610 88.890 ;
        RECT 119.730 85.670 120.250 86.470 ;
        RECT 21.480 82.040 37.140 84.040 ;
        RECT 21.480 78.700 22.940 82.040 ;
        RECT 106.590 81.370 122.250 83.370 ;
        RECT 21.480 76.700 37.140 78.700 ;
        RECT 120.790 78.030 122.250 81.370 ;
        RECT 106.590 76.030 122.250 78.030 ;
        RECT 4.130 60.970 5.780 62.760 ;
        RECT 36.885 53.155 37.405 53.955 ;
        RECT 105.335 53.155 105.855 53.955 ;
        RECT 36.885 48.815 37.405 49.615 ;
        RECT 105.335 48.815 105.855 49.615 ;
        RECT 36.025 46.845 36.405 47.175 ;
        RECT 37.035 46.845 37.415 47.175 ;
        RECT 105.325 46.845 105.705 47.175 ;
        RECT 106.335 46.845 106.715 47.175 ;
        RECT 20.570 44.495 21.200 44.525 ;
        RECT 20.550 43.795 21.200 44.495 ;
        RECT 121.540 44.495 122.170 44.525 ;
        RECT 121.540 43.795 122.190 44.495 ;
        RECT 20.550 43.765 21.180 43.795 ;
        RECT 121.560 43.765 122.190 43.795 ;
        RECT 23.140 42.550 23.520 42.880 ;
        RECT 24.150 42.550 24.530 42.880 ;
        RECT 118.210 42.550 118.590 42.880 ;
        RECT 119.220 42.550 119.600 42.880 ;
        RECT 23.150 40.110 23.670 40.910 ;
        RECT 119.070 40.110 119.590 40.910 ;
        RECT 28.790 36.990 36.960 38.990 ;
        RECT 105.780 36.990 113.950 38.990 ;
        RECT 23.150 35.770 23.670 36.570 ;
        RECT 119.070 35.770 119.590 36.570 ;
        RECT 21.150 31.470 36.810 33.470 ;
        RECT 105.930 31.470 121.590 33.470 ;
        RECT 21.150 28.130 22.610 31.470 ;
        RECT 120.130 28.130 121.590 31.470 ;
        RECT 21.150 26.130 36.810 28.130 ;
        RECT 105.930 26.130 121.590 28.130 ;
      LAYER met3 ;
        RECT 36.175 201.525 37.375 202.325 ;
        RECT 105.695 201.525 106.895 202.325 ;
        RECT 36.175 197.185 37.375 197.985 ;
        RECT 105.695 197.185 106.895 197.985 ;
        RECT 35.715 195.205 37.375 195.555 ;
        RECT 105.695 195.205 107.355 195.555 ;
        RECT 4.110 191.795 5.720 193.165 ;
        RECT 22.990 193.055 37.480 193.065 ;
        RECT 20.170 192.225 37.480 193.055 ;
        RECT 20.170 192.195 24.820 192.225 ;
        RECT 20.170 191.975 24.140 192.195 ;
        RECT 25.860 192.085 37.480 192.225 ;
        RECT 21.910 191.945 24.140 191.975 ;
        RECT 22.460 191.925 24.140 191.945 ;
        RECT 25.910 191.925 37.480 192.085 ;
        RECT 105.590 193.055 120.080 193.065 ;
        RECT 105.590 192.225 122.900 193.055 ;
        RECT 105.590 192.085 117.210 192.225 ;
        RECT 118.250 192.195 122.900 192.225 ;
        RECT 105.590 191.925 117.160 192.085 ;
        RECT 118.930 191.975 122.900 192.195 ;
        RECT 118.930 191.945 121.160 191.975 ;
        RECT 118.930 191.925 120.610 191.945 ;
        RECT 25.910 191.915 27.200 191.925 ;
        RECT 115.870 191.915 117.160 191.925 ;
        RECT 25.910 191.855 26.680 191.915 ;
        RECT 22.520 190.910 24.180 191.260 ;
        RECT 25.920 190.675 26.680 191.855 ;
        RECT 25.850 190.615 26.680 190.675 ;
        RECT 22.520 188.480 23.720 189.280 ;
        RECT 25.550 187.455 26.680 190.615 ;
        RECT 25.620 185.975 26.680 187.455 ;
        RECT 116.390 191.855 117.160 191.915 ;
        RECT 116.390 190.675 117.150 191.855 ;
        RECT 118.890 190.910 120.550 191.260 ;
        RECT 116.390 190.615 117.220 190.675 ;
        RECT 116.390 187.455 117.520 190.615 ;
        RECT 119.350 188.480 120.550 189.280 ;
        RECT 22.520 184.140 23.720 184.940 ;
        RECT 25.550 184.005 26.680 185.975 ;
        RECT 28.460 185.360 35.880 187.360 ;
        RECT 107.190 185.360 114.610 187.360 ;
        RECT 116.390 185.975 117.450 187.455 ;
        RECT 25.370 183.955 27.910 184.005 ;
        RECT 29.020 183.965 31.020 185.360 ;
        RECT 25.370 183.945 28.090 183.955 ;
        RECT 28.580 183.945 31.020 183.965 ;
        RECT 25.370 183.395 31.020 183.945 ;
        RECT 25.550 183.365 31.020 183.395 ;
        RECT 25.550 183.345 28.090 183.365 ;
        RECT 28.580 183.285 31.020 183.365 ;
        RECT 29.020 181.840 31.020 183.285 ;
        RECT 112.050 183.965 114.050 185.360 ;
        RECT 116.390 184.005 117.520 185.975 ;
        RECT 119.350 184.140 120.550 184.940 ;
        RECT 112.050 183.945 114.490 183.965 ;
        RECT 115.160 183.955 117.700 184.005 ;
        RECT 114.980 183.945 117.700 183.955 ;
        RECT 112.050 183.395 117.700 183.945 ;
        RECT 112.050 183.365 117.520 183.395 ;
        RECT 112.050 183.285 114.490 183.365 ;
        RECT 114.980 183.345 117.520 183.365 ;
        RECT 112.050 181.840 114.050 183.285 ;
        RECT 20.820 179.840 36.480 181.840 ;
        RECT 106.590 179.840 122.250 181.840 ;
        RECT 4.130 171.350 5.780 173.140 ;
        RECT 36.175 151.955 37.375 152.755 ;
        RECT 105.695 151.955 106.895 152.755 ;
        RECT 36.175 147.615 37.375 148.415 ;
        RECT 105.695 147.615 106.895 148.415 ;
        RECT 35.715 145.635 37.375 145.985 ;
        RECT 105.695 145.635 107.355 145.985 ;
        RECT 22.990 143.485 37.480 143.495 ;
        RECT 20.170 142.655 37.480 143.485 ;
        RECT 20.170 142.625 24.820 142.655 ;
        RECT 20.170 142.405 24.140 142.625 ;
        RECT 25.860 142.515 37.480 142.655 ;
        RECT 21.910 142.375 24.140 142.405 ;
        RECT 22.460 142.355 24.140 142.375 ;
        RECT 25.910 142.355 37.480 142.515 ;
        RECT 105.590 143.485 120.080 143.495 ;
        RECT 105.590 142.655 122.900 143.485 ;
        RECT 105.590 142.515 117.210 142.655 ;
        RECT 118.250 142.625 122.900 142.655 ;
        RECT 105.590 142.355 117.160 142.515 ;
        RECT 118.930 142.405 122.900 142.625 ;
        RECT 118.930 142.375 121.160 142.405 ;
        RECT 118.930 142.355 120.610 142.375 ;
        RECT 25.910 142.345 27.200 142.355 ;
        RECT 115.870 142.345 117.160 142.355 ;
        RECT 25.910 142.285 26.680 142.345 ;
        RECT 22.520 141.340 24.180 141.690 ;
        RECT 25.920 141.105 26.680 142.285 ;
        RECT 25.850 141.045 26.680 141.105 ;
        RECT 22.520 138.910 23.720 139.710 ;
        RECT 25.550 137.885 26.680 141.045 ;
        RECT 25.620 136.405 26.680 137.885 ;
        RECT 116.390 142.285 117.160 142.345 ;
        RECT 116.390 141.105 117.150 142.285 ;
        RECT 118.890 141.340 120.550 141.690 ;
        RECT 116.390 141.045 117.220 141.105 ;
        RECT 116.390 137.885 117.520 141.045 ;
        RECT 119.350 138.910 120.550 139.710 ;
        RECT 22.520 134.570 23.720 135.370 ;
        RECT 25.550 134.435 26.680 136.405 ;
        RECT 28.460 135.790 35.880 137.790 ;
        RECT 107.190 135.790 114.610 137.790 ;
        RECT 116.390 136.405 117.450 137.885 ;
        RECT 25.370 134.385 27.910 134.435 ;
        RECT 29.020 134.395 31.020 135.790 ;
        RECT 25.370 134.375 28.090 134.385 ;
        RECT 28.580 134.375 31.020 134.395 ;
        RECT 25.370 133.825 31.020 134.375 ;
        RECT 25.550 133.795 31.020 133.825 ;
        RECT 25.550 133.775 28.090 133.795 ;
        RECT 28.580 133.715 31.020 133.795 ;
        RECT 29.020 132.270 31.020 133.715 ;
        RECT 112.050 134.395 114.050 135.790 ;
        RECT 116.390 134.435 117.520 136.405 ;
        RECT 119.350 134.570 120.550 135.370 ;
        RECT 112.050 134.375 114.490 134.395 ;
        RECT 115.160 134.385 117.700 134.435 ;
        RECT 114.980 134.375 117.700 134.385 ;
        RECT 112.050 133.825 117.700 134.375 ;
        RECT 112.050 133.795 117.520 133.825 ;
        RECT 112.050 133.715 114.490 133.795 ;
        RECT 114.980 133.775 117.520 133.795 ;
        RECT 112.050 132.270 114.050 133.715 ;
        RECT 20.820 130.270 36.480 132.270 ;
        RECT 106.590 130.270 122.250 132.270 ;
        RECT 4.160 113.000 5.810 114.790 ;
        RECT 36.835 103.725 38.035 104.525 ;
        RECT 105.695 103.055 106.895 103.855 ;
        RECT 36.835 99.385 38.035 100.185 ;
        RECT 105.695 98.715 106.895 99.515 ;
        RECT 36.375 97.405 38.035 97.755 ;
        RECT 105.695 96.735 107.355 97.085 ;
        RECT 23.650 95.255 38.140 95.265 ;
        RECT 20.830 94.425 38.140 95.255 ;
        RECT 20.830 94.395 25.480 94.425 ;
        RECT 20.830 94.175 24.800 94.395 ;
        RECT 26.520 94.285 38.140 94.425 ;
        RECT 22.570 94.145 24.800 94.175 ;
        RECT 23.120 94.125 24.800 94.145 ;
        RECT 26.570 94.125 38.140 94.285 ;
        RECT 105.590 94.585 120.080 94.595 ;
        RECT 26.570 94.115 27.860 94.125 ;
        RECT 26.570 94.055 27.340 94.115 ;
        RECT 23.180 93.110 24.840 93.460 ;
        RECT 26.580 92.875 27.340 94.055 ;
        RECT 105.590 93.755 122.900 94.585 ;
        RECT 105.590 93.615 117.210 93.755 ;
        RECT 118.250 93.725 122.900 93.755 ;
        RECT 105.590 93.455 117.160 93.615 ;
        RECT 118.930 93.505 122.900 93.725 ;
        RECT 118.930 93.475 121.160 93.505 ;
        RECT 118.930 93.455 120.610 93.475 ;
        RECT 115.870 93.445 117.160 93.455 ;
        RECT 26.510 92.815 27.340 92.875 ;
        RECT 23.180 90.680 24.380 91.480 ;
        RECT 26.210 89.655 27.340 92.815 ;
        RECT 26.280 88.175 27.340 89.655 ;
        RECT 116.390 93.385 117.160 93.445 ;
        RECT 116.390 92.205 117.150 93.385 ;
        RECT 118.890 92.440 120.550 92.790 ;
        RECT 116.390 92.145 117.220 92.205 ;
        RECT 23.180 86.340 24.380 87.140 ;
        RECT 26.210 86.205 27.340 88.175 ;
        RECT 29.120 87.560 36.540 89.560 ;
        RECT 116.390 88.985 117.520 92.145 ;
        RECT 119.350 90.010 120.550 90.810 ;
        RECT 26.030 86.155 28.570 86.205 ;
        RECT 29.680 86.165 31.680 87.560 ;
        RECT 107.190 86.890 114.610 88.890 ;
        RECT 116.390 87.505 117.450 88.985 ;
        RECT 26.030 86.145 28.750 86.155 ;
        RECT 29.240 86.145 31.680 86.165 ;
        RECT 26.030 85.595 31.680 86.145 ;
        RECT 26.210 85.565 31.680 85.595 ;
        RECT 26.210 85.545 28.750 85.565 ;
        RECT 29.240 85.485 31.680 85.565 ;
        RECT 29.680 84.040 31.680 85.485 ;
        RECT 112.050 85.495 114.050 86.890 ;
        RECT 116.390 85.535 117.520 87.505 ;
        RECT 119.350 85.670 120.550 86.470 ;
        RECT 112.050 85.475 114.490 85.495 ;
        RECT 115.160 85.485 117.700 85.535 ;
        RECT 114.980 85.475 117.700 85.485 ;
        RECT 112.050 84.925 117.700 85.475 ;
        RECT 112.050 84.895 117.520 84.925 ;
        RECT 112.050 84.815 114.490 84.895 ;
        RECT 114.980 84.875 117.520 84.895 ;
        RECT 21.480 82.040 37.140 84.040 ;
        RECT 112.050 83.370 114.050 84.815 ;
        RECT 106.590 81.370 122.250 83.370 ;
        RECT 4.130 60.970 5.780 62.760 ;
        RECT 36.505 53.155 37.705 53.955 ;
        RECT 105.035 53.155 106.235 53.955 ;
        RECT 36.505 48.815 37.705 49.615 ;
        RECT 105.035 48.815 106.235 49.615 ;
        RECT 36.045 46.835 37.705 47.185 ;
        RECT 105.035 46.835 106.695 47.185 ;
        RECT 23.320 44.685 37.810 44.695 ;
        RECT 20.500 43.855 37.810 44.685 ;
        RECT 20.500 43.825 25.150 43.855 ;
        RECT 20.500 43.605 24.470 43.825 ;
        RECT 26.190 43.715 37.810 43.855 ;
        RECT 22.240 43.575 24.470 43.605 ;
        RECT 22.790 43.555 24.470 43.575 ;
        RECT 26.240 43.555 37.810 43.715 ;
        RECT 104.930 44.685 119.420 44.695 ;
        RECT 104.930 43.855 122.240 44.685 ;
        RECT 104.930 43.715 116.550 43.855 ;
        RECT 117.590 43.825 122.240 43.855 ;
        RECT 104.930 43.555 116.500 43.715 ;
        RECT 118.270 43.605 122.240 43.825 ;
        RECT 118.270 43.575 120.500 43.605 ;
        RECT 118.270 43.555 119.950 43.575 ;
        RECT 26.240 43.545 27.530 43.555 ;
        RECT 115.210 43.545 116.500 43.555 ;
        RECT 26.240 43.485 27.010 43.545 ;
        RECT 22.850 42.540 24.510 42.890 ;
        RECT 26.250 42.305 27.010 43.485 ;
        RECT 26.180 42.245 27.010 42.305 ;
        RECT 22.850 40.110 24.050 40.910 ;
        RECT 25.880 39.085 27.010 42.245 ;
        RECT 25.950 37.605 27.010 39.085 ;
        RECT 115.730 43.485 116.500 43.545 ;
        RECT 115.730 42.305 116.490 43.485 ;
        RECT 118.230 42.540 119.890 42.890 ;
        RECT 115.730 42.245 116.560 42.305 ;
        RECT 115.730 39.085 116.860 42.245 ;
        RECT 118.690 40.110 119.890 40.910 ;
        RECT 22.850 35.770 24.050 36.570 ;
        RECT 25.880 35.635 27.010 37.605 ;
        RECT 28.790 36.990 36.210 38.990 ;
        RECT 106.530 36.990 113.950 38.990 ;
        RECT 115.730 37.605 116.790 39.085 ;
        RECT 25.700 35.585 28.240 35.635 ;
        RECT 29.350 35.595 31.350 36.990 ;
        RECT 25.700 35.575 28.420 35.585 ;
        RECT 28.910 35.575 31.350 35.595 ;
        RECT 25.700 35.025 31.350 35.575 ;
        RECT 25.880 34.995 31.350 35.025 ;
        RECT 25.880 34.975 28.420 34.995 ;
        RECT 28.910 34.915 31.350 34.995 ;
        RECT 29.350 33.470 31.350 34.915 ;
        RECT 111.390 35.595 113.390 36.990 ;
        RECT 115.730 35.635 116.860 37.605 ;
        RECT 118.690 35.770 119.890 36.570 ;
        RECT 111.390 35.575 113.830 35.595 ;
        RECT 114.500 35.585 117.040 35.635 ;
        RECT 114.320 35.575 117.040 35.585 ;
        RECT 111.390 35.025 117.040 35.575 ;
        RECT 111.390 34.995 116.860 35.025 ;
        RECT 111.390 34.915 113.830 34.995 ;
        RECT 114.320 34.975 116.860 34.995 ;
        RECT 111.390 33.470 113.390 34.915 ;
        RECT 21.150 31.470 36.810 33.470 ;
        RECT 105.930 31.470 121.590 33.470 ;
      LAYER met4 ;
        RECT 4.000 115.400 6.000 220.760 ;
        RECT 36.175 194.835 37.375 216.365 ;
        RECT 105.695 194.835 106.895 216.365 ;
        RECT 36.175 194.625 37.380 194.835 ;
        RECT 22.500 191.860 23.690 193.055 ;
        RECT 36.170 192.115 37.380 194.625 ;
        RECT 105.690 194.625 106.895 194.835 ;
        RECT 105.690 192.115 106.900 194.625 ;
        RECT 36.170 191.905 37.370 192.115 ;
        RECT 105.700 191.905 106.900 192.115 ;
        RECT 119.380 191.860 120.570 193.055 ;
        RECT 22.500 191.825 23.720 191.860 ;
        RECT 22.520 170.100 23.720 191.825 ;
        RECT 119.350 191.825 120.570 191.860 ;
        RECT 29.570 181.860 30.470 183.860 ;
        RECT 112.600 181.860 113.500 183.860 ;
        RECT 119.350 170.100 120.550 191.825 ;
        RECT 36.175 145.265 37.375 166.795 ;
        RECT 105.695 145.265 106.895 166.795 ;
        RECT 36.175 145.055 37.380 145.265 ;
        RECT 22.500 142.290 23.690 143.485 ;
        RECT 36.170 142.545 37.380 145.055 ;
        RECT 105.690 145.055 106.895 145.265 ;
        RECT 105.690 142.545 106.900 145.055 ;
        RECT 36.170 142.335 37.370 142.545 ;
        RECT 105.700 142.335 106.900 142.545 ;
        RECT 119.380 142.290 120.570 143.485 ;
        RECT 22.500 142.255 23.720 142.290 ;
        RECT 22.520 120.530 23.720 142.255 ;
        RECT 119.350 142.255 120.570 142.290 ;
        RECT 29.570 132.290 30.470 134.290 ;
        RECT 112.600 132.290 113.500 134.290 ;
        RECT 119.350 120.530 120.550 142.255 ;
        RECT 4.000 112.600 6.030 115.400 ;
        RECT 4.000 103.450 6.000 112.600 ;
        RECT 4.000 101.970 6.050 103.450 ;
        RECT 4.000 69.170 6.000 101.970 ;
        RECT 36.835 97.035 38.035 118.565 ;
        RECT 36.835 96.825 38.040 97.035 ;
        RECT 23.160 94.060 24.350 95.255 ;
        RECT 36.830 94.315 38.040 96.825 ;
        RECT 105.695 96.365 106.895 117.895 ;
        RECT 105.690 96.155 106.895 96.365 ;
        RECT 36.830 94.105 38.030 94.315 ;
        RECT 23.160 94.025 24.380 94.060 ;
        RECT 23.180 72.300 24.380 94.025 ;
        RECT 105.690 93.645 106.900 96.155 ;
        RECT 105.700 93.435 106.900 93.645 ;
        RECT 119.380 93.390 120.570 94.585 ;
        RECT 119.350 93.355 120.570 93.390 ;
        RECT 30.230 84.060 31.130 86.060 ;
        RECT 112.600 83.390 113.500 85.390 ;
        RECT 119.350 71.630 120.550 93.355 ;
        RECT 4.000 67.690 6.010 69.170 ;
        RECT 4.000 5.000 6.000 67.690 ;
        RECT 36.505 46.465 37.705 67.995 ;
        RECT 105.035 46.465 106.235 67.995 ;
        RECT 36.505 46.255 37.710 46.465 ;
        RECT 22.830 43.490 24.020 44.685 ;
        RECT 36.500 43.745 37.710 46.255 ;
        RECT 105.030 46.255 106.235 46.465 ;
        RECT 105.030 43.745 106.240 46.255 ;
        RECT 36.500 43.535 37.700 43.745 ;
        RECT 105.040 43.535 106.240 43.745 ;
        RECT 118.720 43.490 119.910 44.685 ;
        RECT 22.830 43.455 24.050 43.490 ;
        RECT 22.850 21.730 24.050 43.455 ;
        RECT 118.690 43.455 119.910 43.490 ;
        RECT 29.900 33.490 30.800 35.490 ;
        RECT 111.940 33.490 112.840 35.490 ;
        RECT 118.690 21.730 119.890 43.455 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 21.615 203.145 38.125 216.115 ;
        RECT 104.945 203.145 121.455 216.115 ;
        RECT 34.665 198.365 38.695 201.145 ;
        RECT 104.375 198.365 108.405 201.145 ;
        RECT 21.200 185.320 25.230 188.100 ;
        RECT 117.840 185.320 121.870 188.100 ;
        RECT 21.770 170.350 38.280 183.320 ;
        RECT 104.790 170.350 121.300 183.320 ;
        RECT 21.615 153.575 38.125 166.545 ;
        RECT 104.945 153.575 121.455 166.545 ;
        RECT 34.665 148.795 38.695 151.575 ;
        RECT 104.375 148.795 108.405 151.575 ;
        RECT 21.200 135.750 25.230 138.530 ;
        RECT 117.840 135.750 121.870 138.530 ;
        RECT 21.770 120.780 38.280 133.750 ;
        RECT 104.790 120.780 121.300 133.750 ;
        RECT 22.275 105.345 38.785 118.315 ;
        RECT 104.945 104.675 121.455 117.645 ;
        RECT 35.325 100.565 39.355 103.345 ;
        RECT 104.375 99.895 108.405 102.675 ;
        RECT 21.860 87.520 25.890 90.300 ;
        RECT 117.840 86.850 121.870 89.630 ;
        RECT 22.430 72.550 38.940 85.520 ;
        RECT 104.790 71.880 121.300 84.850 ;
        RECT 21.945 54.775 38.455 67.745 ;
        RECT 104.285 54.775 120.795 67.745 ;
        RECT 34.995 49.995 39.025 52.775 ;
        RECT 103.715 49.995 107.745 52.775 ;
        RECT 21.530 36.950 25.560 39.730 ;
        RECT 117.180 36.950 121.210 39.730 ;
        RECT 22.100 21.980 38.610 34.950 ;
        RECT 104.130 21.980 120.640 34.950 ;
      LAYER li1 ;
        RECT 22.005 215.555 37.735 215.725 ;
        RECT 22.005 203.705 22.175 215.555 ;
        RECT 23.465 204.610 23.635 214.650 ;
        RECT 25.045 204.610 25.215 214.650 ;
        RECT 26.625 204.610 26.795 214.650 ;
        RECT 28.205 204.610 28.375 214.650 ;
        RECT 29.785 204.610 29.955 214.650 ;
        RECT 31.365 204.610 31.535 214.650 ;
        RECT 32.945 204.610 33.115 214.650 ;
        RECT 34.525 204.610 34.695 214.650 ;
        RECT 36.105 204.610 36.275 214.650 ;
        RECT 37.565 203.705 37.735 215.555 ;
        RECT 22.005 203.535 37.735 203.705 ;
        RECT 105.335 215.555 121.065 215.725 ;
        RECT 105.335 203.705 105.505 215.555 ;
        RECT 106.795 204.610 106.965 214.650 ;
        RECT 108.375 204.610 108.545 214.650 ;
        RECT 109.955 204.610 110.125 214.650 ;
        RECT 111.535 204.610 111.705 214.650 ;
        RECT 113.115 204.610 113.285 214.650 ;
        RECT 114.695 204.610 114.865 214.650 ;
        RECT 116.275 204.610 116.445 214.650 ;
        RECT 117.855 204.610 118.025 214.650 ;
        RECT 119.435 204.610 119.605 214.650 ;
        RECT 120.895 203.705 121.065 215.555 ;
        RECT 105.335 203.535 121.065 203.705 ;
        RECT 23.315 196.085 23.485 201.125 ;
        RECT 24.895 196.085 25.065 201.125 ;
        RECT 26.475 196.085 26.645 201.125 ;
        RECT 28.055 196.085 28.225 201.125 ;
        RECT 29.635 196.085 29.805 201.125 ;
        RECT 31.215 196.085 31.385 201.125 ;
        RECT 35.055 200.085 35.225 200.855 ;
        RECT 36.635 200.085 36.805 200.855 ;
        RECT 106.265 200.085 106.435 200.855 ;
        RECT 107.845 200.085 108.015 200.855 ;
        RECT 35.035 199.425 37.275 200.085 ;
        RECT 105.795 199.425 108.035 200.085 ;
        RECT 35.055 198.655 35.225 199.425 ;
        RECT 36.635 198.655 36.805 199.425 ;
        RECT 106.265 198.655 106.435 199.425 ;
        RECT 107.845 198.655 108.015 199.425 ;
        RECT 111.685 196.085 111.855 201.125 ;
        RECT 113.265 196.085 113.435 201.125 ;
        RECT 114.845 196.085 115.015 201.125 ;
        RECT 116.425 196.085 116.595 201.125 ;
        RECT 118.005 196.085 118.175 201.125 ;
        RECT 119.585 196.085 119.755 201.125 ;
        RECT 23.090 187.040 23.260 187.810 ;
        RECT 24.670 187.040 24.840 187.810 ;
        RECT 118.230 187.040 118.400 187.810 ;
        RECT 119.810 187.040 119.980 187.810 ;
        RECT 22.620 186.380 24.860 187.040 ;
        RECT 118.210 186.380 120.450 187.040 ;
        RECT 23.090 185.610 23.260 186.380 ;
        RECT 24.670 185.610 24.840 186.380 ;
        RECT 118.230 185.610 118.400 186.380 ;
        RECT 119.810 185.610 119.980 186.380 ;
        RECT 22.160 182.760 37.890 182.930 ;
        RECT 22.160 170.910 22.330 182.760 ;
        RECT 37.720 170.910 37.890 182.760 ;
        RECT 22.160 170.740 37.890 170.910 ;
        RECT 105.180 182.760 120.910 182.930 ;
        RECT 105.180 170.910 105.350 182.760 ;
        RECT 120.740 170.910 120.910 182.760 ;
        RECT 105.180 170.740 120.910 170.910 ;
        RECT 22.005 165.985 37.735 166.155 ;
        RECT 22.005 154.135 22.175 165.985 ;
        RECT 23.465 155.040 23.635 165.080 ;
        RECT 25.045 155.040 25.215 165.080 ;
        RECT 26.625 155.040 26.795 165.080 ;
        RECT 28.205 155.040 28.375 165.080 ;
        RECT 29.785 155.040 29.955 165.080 ;
        RECT 31.365 155.040 31.535 165.080 ;
        RECT 32.945 155.040 33.115 165.080 ;
        RECT 34.525 155.040 34.695 165.080 ;
        RECT 36.105 155.040 36.275 165.080 ;
        RECT 37.565 154.135 37.735 165.985 ;
        RECT 22.005 153.965 37.735 154.135 ;
        RECT 105.335 165.985 121.065 166.155 ;
        RECT 105.335 154.135 105.505 165.985 ;
        RECT 106.795 155.040 106.965 165.080 ;
        RECT 108.375 155.040 108.545 165.080 ;
        RECT 109.955 155.040 110.125 165.080 ;
        RECT 111.535 155.040 111.705 165.080 ;
        RECT 113.115 155.040 113.285 165.080 ;
        RECT 114.695 155.040 114.865 165.080 ;
        RECT 116.275 155.040 116.445 165.080 ;
        RECT 117.855 155.040 118.025 165.080 ;
        RECT 119.435 155.040 119.605 165.080 ;
        RECT 120.895 154.135 121.065 165.985 ;
        RECT 105.335 153.965 121.065 154.135 ;
        RECT 23.315 146.515 23.485 151.555 ;
        RECT 24.895 146.515 25.065 151.555 ;
        RECT 26.475 146.515 26.645 151.555 ;
        RECT 28.055 146.515 28.225 151.555 ;
        RECT 29.635 146.515 29.805 151.555 ;
        RECT 31.215 146.515 31.385 151.555 ;
        RECT 35.055 150.515 35.225 151.285 ;
        RECT 36.635 150.515 36.805 151.285 ;
        RECT 106.265 150.515 106.435 151.285 ;
        RECT 107.845 150.515 108.015 151.285 ;
        RECT 35.035 149.855 37.275 150.515 ;
        RECT 105.795 149.855 108.035 150.515 ;
        RECT 35.055 149.085 35.225 149.855 ;
        RECT 36.635 149.085 36.805 149.855 ;
        RECT 106.265 149.085 106.435 149.855 ;
        RECT 107.845 149.085 108.015 149.855 ;
        RECT 111.685 146.515 111.855 151.555 ;
        RECT 113.265 146.515 113.435 151.555 ;
        RECT 114.845 146.515 115.015 151.555 ;
        RECT 116.425 146.515 116.595 151.555 ;
        RECT 118.005 146.515 118.175 151.555 ;
        RECT 119.585 146.515 119.755 151.555 ;
        RECT 23.090 137.470 23.260 138.240 ;
        RECT 24.670 137.470 24.840 138.240 ;
        RECT 118.230 137.470 118.400 138.240 ;
        RECT 119.810 137.470 119.980 138.240 ;
        RECT 22.620 136.810 24.860 137.470 ;
        RECT 118.210 136.810 120.450 137.470 ;
        RECT 23.090 136.040 23.260 136.810 ;
        RECT 24.670 136.040 24.840 136.810 ;
        RECT 118.230 136.040 118.400 136.810 ;
        RECT 119.810 136.040 119.980 136.810 ;
        RECT 22.160 133.190 37.890 133.360 ;
        RECT 22.160 121.340 22.330 133.190 ;
        RECT 37.720 121.340 37.890 133.190 ;
        RECT 22.160 121.170 37.890 121.340 ;
        RECT 105.180 133.190 120.910 133.360 ;
        RECT 105.180 121.340 105.350 133.190 ;
        RECT 120.740 121.340 120.910 133.190 ;
        RECT 105.180 121.170 120.910 121.340 ;
        RECT 22.665 117.755 38.395 117.925 ;
        RECT 22.665 105.905 22.835 117.755 ;
        RECT 24.125 106.810 24.295 116.850 ;
        RECT 25.705 106.810 25.875 116.850 ;
        RECT 27.285 106.810 27.455 116.850 ;
        RECT 28.865 106.810 29.035 116.850 ;
        RECT 30.445 106.810 30.615 116.850 ;
        RECT 32.025 106.810 32.195 116.850 ;
        RECT 33.605 106.810 33.775 116.850 ;
        RECT 35.185 106.810 35.355 116.850 ;
        RECT 36.765 106.810 36.935 116.850 ;
        RECT 38.225 105.905 38.395 117.755 ;
        RECT 22.665 105.735 38.395 105.905 ;
        RECT 105.335 117.085 121.065 117.255 ;
        RECT 105.335 105.235 105.505 117.085 ;
        RECT 106.795 106.140 106.965 116.180 ;
        RECT 108.375 106.140 108.545 116.180 ;
        RECT 109.955 106.140 110.125 116.180 ;
        RECT 111.535 106.140 111.705 116.180 ;
        RECT 113.115 106.140 113.285 116.180 ;
        RECT 114.695 106.140 114.865 116.180 ;
        RECT 116.275 106.140 116.445 116.180 ;
        RECT 117.855 106.140 118.025 116.180 ;
        RECT 119.435 106.140 119.605 116.180 ;
        RECT 120.895 105.235 121.065 117.085 ;
        RECT 105.335 105.065 121.065 105.235 ;
        RECT 23.975 98.285 24.145 103.325 ;
        RECT 25.555 98.285 25.725 103.325 ;
        RECT 27.135 98.285 27.305 103.325 ;
        RECT 28.715 98.285 28.885 103.325 ;
        RECT 30.295 98.285 30.465 103.325 ;
        RECT 31.875 98.285 32.045 103.325 ;
        RECT 35.715 102.285 35.885 103.055 ;
        RECT 37.295 102.285 37.465 103.055 ;
        RECT 35.695 101.625 37.935 102.285 ;
        RECT 35.715 100.855 35.885 101.625 ;
        RECT 37.295 100.855 37.465 101.625 ;
        RECT 106.265 101.615 106.435 102.385 ;
        RECT 107.845 101.615 108.015 102.385 ;
        RECT 105.795 100.955 108.035 101.615 ;
        RECT 106.265 100.185 106.435 100.955 ;
        RECT 107.845 100.185 108.015 100.955 ;
        RECT 111.685 97.615 111.855 102.655 ;
        RECT 113.265 97.615 113.435 102.655 ;
        RECT 114.845 97.615 115.015 102.655 ;
        RECT 116.425 97.615 116.595 102.655 ;
        RECT 118.005 97.615 118.175 102.655 ;
        RECT 119.585 97.615 119.755 102.655 ;
        RECT 23.750 89.240 23.920 90.010 ;
        RECT 25.330 89.240 25.500 90.010 ;
        RECT 23.280 88.580 25.520 89.240 ;
        RECT 23.750 87.810 23.920 88.580 ;
        RECT 25.330 87.810 25.500 88.580 ;
        RECT 118.230 88.570 118.400 89.340 ;
        RECT 119.810 88.570 119.980 89.340 ;
        RECT 118.210 87.910 120.450 88.570 ;
        RECT 118.230 87.140 118.400 87.910 ;
        RECT 119.810 87.140 119.980 87.910 ;
        RECT 22.820 84.960 38.550 85.130 ;
        RECT 22.820 73.110 22.990 84.960 ;
        RECT 38.380 73.110 38.550 84.960 ;
        RECT 22.820 72.940 38.550 73.110 ;
        RECT 105.180 84.290 120.910 84.460 ;
        RECT 105.180 72.440 105.350 84.290 ;
        RECT 120.740 72.440 120.910 84.290 ;
        RECT 105.180 72.270 120.910 72.440 ;
        RECT 22.335 67.185 38.065 67.355 ;
        RECT 22.335 55.335 22.505 67.185 ;
        RECT 23.795 56.240 23.965 66.280 ;
        RECT 25.375 56.240 25.545 66.280 ;
        RECT 26.955 56.240 27.125 66.280 ;
        RECT 28.535 56.240 28.705 66.280 ;
        RECT 30.115 56.240 30.285 66.280 ;
        RECT 31.695 56.240 31.865 66.280 ;
        RECT 33.275 56.240 33.445 66.280 ;
        RECT 34.855 56.240 35.025 66.280 ;
        RECT 36.435 56.240 36.605 66.280 ;
        RECT 37.895 55.335 38.065 67.185 ;
        RECT 22.335 55.165 38.065 55.335 ;
        RECT 104.675 67.185 120.405 67.355 ;
        RECT 104.675 55.335 104.845 67.185 ;
        RECT 106.135 56.240 106.305 66.280 ;
        RECT 107.715 56.240 107.885 66.280 ;
        RECT 109.295 56.240 109.465 66.280 ;
        RECT 110.875 56.240 111.045 66.280 ;
        RECT 112.455 56.240 112.625 66.280 ;
        RECT 114.035 56.240 114.205 66.280 ;
        RECT 115.615 56.240 115.785 66.280 ;
        RECT 117.195 56.240 117.365 66.280 ;
        RECT 118.775 56.240 118.945 66.280 ;
        RECT 120.235 55.335 120.405 67.185 ;
        RECT 104.675 55.165 120.405 55.335 ;
        RECT 23.645 47.715 23.815 52.755 ;
        RECT 25.225 47.715 25.395 52.755 ;
        RECT 26.805 47.715 26.975 52.755 ;
        RECT 28.385 47.715 28.555 52.755 ;
        RECT 29.965 47.715 30.135 52.755 ;
        RECT 31.545 47.715 31.715 52.755 ;
        RECT 35.385 51.715 35.555 52.485 ;
        RECT 36.965 51.715 37.135 52.485 ;
        RECT 105.605 51.715 105.775 52.485 ;
        RECT 107.185 51.715 107.355 52.485 ;
        RECT 35.365 51.055 37.605 51.715 ;
        RECT 105.135 51.055 107.375 51.715 ;
        RECT 35.385 50.285 35.555 51.055 ;
        RECT 36.965 50.285 37.135 51.055 ;
        RECT 105.605 50.285 105.775 51.055 ;
        RECT 107.185 50.285 107.355 51.055 ;
        RECT 111.025 47.715 111.195 52.755 ;
        RECT 112.605 47.715 112.775 52.755 ;
        RECT 114.185 47.715 114.355 52.755 ;
        RECT 115.765 47.715 115.935 52.755 ;
        RECT 117.345 47.715 117.515 52.755 ;
        RECT 118.925 47.715 119.095 52.755 ;
        RECT 23.420 38.670 23.590 39.440 ;
        RECT 25.000 38.670 25.170 39.440 ;
        RECT 117.570 38.670 117.740 39.440 ;
        RECT 119.150 38.670 119.320 39.440 ;
        RECT 22.950 38.010 25.190 38.670 ;
        RECT 117.550 38.010 119.790 38.670 ;
        RECT 23.420 37.240 23.590 38.010 ;
        RECT 25.000 37.240 25.170 38.010 ;
        RECT 117.570 37.240 117.740 38.010 ;
        RECT 119.150 37.240 119.320 38.010 ;
        RECT 22.490 34.390 38.220 34.560 ;
        RECT 22.490 22.540 22.660 34.390 ;
        RECT 38.050 22.540 38.220 34.390 ;
        RECT 22.490 22.370 38.220 22.540 ;
        RECT 104.520 34.390 120.250 34.560 ;
        RECT 104.520 22.540 104.690 34.390 ;
        RECT 120.080 22.540 120.250 34.390 ;
        RECT 104.520 22.370 120.250 22.540 ;
      LAYER met1 ;
        RECT 21.945 215.525 37.795 215.755 ;
        RECT 105.275 215.525 121.125 215.755 ;
        RECT 21.945 203.735 22.235 215.525 ;
        RECT 23.415 204.625 23.685 214.635 ;
        RECT 24.995 204.625 25.265 214.635 ;
        RECT 26.575 204.625 26.845 214.635 ;
        RECT 28.155 204.625 28.425 214.635 ;
        RECT 29.735 204.625 30.005 214.635 ;
        RECT 31.315 204.625 31.585 214.635 ;
        RECT 32.895 204.625 33.165 214.635 ;
        RECT 34.475 204.625 34.745 214.635 ;
        RECT 36.055 204.625 36.325 214.635 ;
        RECT 106.745 204.625 107.015 214.635 ;
        RECT 108.325 204.625 108.595 214.635 ;
        RECT 109.905 204.625 110.175 214.635 ;
        RECT 111.485 204.625 111.755 214.635 ;
        RECT 113.065 204.625 113.335 214.635 ;
        RECT 114.645 204.625 114.915 214.635 ;
        RECT 116.225 204.625 116.495 214.635 ;
        RECT 117.805 204.625 118.075 214.635 ;
        RECT 119.385 204.625 119.655 214.635 ;
        RECT 34.585 203.735 35.765 203.785 ;
        RECT 107.305 203.735 108.485 203.785 ;
        RECT 120.835 203.735 121.125 215.525 ;
        RECT 21.945 203.505 37.795 203.735 ;
        RECT 105.275 203.505 121.125 203.735 ;
        RECT 34.585 203.455 35.765 203.505 ;
        RECT 107.305 203.455 108.485 203.505 ;
        RECT 23.265 196.105 23.535 201.105 ;
        RECT 24.845 196.105 25.115 201.105 ;
        RECT 26.425 196.105 26.695 201.105 ;
        RECT 28.005 196.105 28.275 201.105 ;
        RECT 29.585 196.105 29.855 201.105 ;
        RECT 31.165 196.105 31.435 201.105 ;
        RECT 35.025 200.195 35.255 200.855 ;
        RECT 36.605 200.195 36.835 200.855 ;
        RECT 35.025 199.315 36.835 200.195 ;
        RECT 35.025 198.655 35.255 199.315 ;
        RECT 36.605 198.655 36.835 199.315 ;
        RECT 106.235 200.195 106.465 200.855 ;
        RECT 107.815 200.195 108.045 200.855 ;
        RECT 106.235 199.315 108.045 200.195 ;
        RECT 106.235 198.655 106.465 199.315 ;
        RECT 107.815 198.655 108.045 199.315 ;
        RECT 111.635 196.105 111.905 201.105 ;
        RECT 113.215 196.105 113.485 201.105 ;
        RECT 114.795 196.105 115.065 201.105 ;
        RECT 116.375 196.105 116.645 201.105 ;
        RECT 117.955 196.105 118.225 201.105 ;
        RECT 119.535 196.105 119.805 201.105 ;
        RECT 20.750 194.515 21.910 194.535 ;
        RECT 19.590 194.485 21.910 194.515 ;
        RECT 121.160 194.515 122.320 194.535 ;
        RECT 121.160 194.485 123.480 194.515 ;
        RECT 19.590 193.565 22.240 194.485 ;
        RECT 120.830 193.565 123.480 194.485 ;
        RECT 19.590 193.535 21.910 193.565 ;
        RECT 121.160 193.535 123.480 193.565 ;
        RECT 19.590 193.515 21.100 193.535 ;
        RECT 121.970 193.515 123.480 193.535 ;
        RECT 23.060 187.150 23.290 187.810 ;
        RECT 24.640 187.150 24.870 187.810 ;
        RECT 23.060 186.270 24.870 187.150 ;
        RECT 23.060 185.610 23.290 186.270 ;
        RECT 24.640 185.610 24.870 186.270 ;
        RECT 118.200 187.150 118.430 187.810 ;
        RECT 119.780 187.150 120.010 187.810 ;
        RECT 118.200 186.270 120.010 187.150 ;
        RECT 118.200 185.610 118.430 186.270 ;
        RECT 119.780 185.610 120.010 186.270 ;
        RECT 24.130 182.960 25.310 183.010 ;
        RECT 117.760 182.960 118.940 183.010 ;
        RECT 22.100 182.730 37.950 182.960 ;
        RECT 24.130 182.680 25.310 182.730 ;
        RECT 37.660 170.940 37.950 182.730 ;
        RECT 22.100 170.710 37.950 170.940 ;
        RECT 105.120 182.730 120.970 182.960 ;
        RECT 105.120 170.940 105.410 182.730 ;
        RECT 117.760 182.680 118.940 182.730 ;
        RECT 105.120 170.710 120.970 170.940 ;
        RECT 21.945 165.955 37.795 166.185 ;
        RECT 105.275 165.955 121.125 166.185 ;
        RECT 21.945 154.165 22.235 165.955 ;
        RECT 23.415 155.055 23.685 165.065 ;
        RECT 24.995 155.055 25.265 165.065 ;
        RECT 26.575 155.055 26.845 165.065 ;
        RECT 28.155 155.055 28.425 165.065 ;
        RECT 29.735 155.055 30.005 165.065 ;
        RECT 31.315 155.055 31.585 165.065 ;
        RECT 32.895 155.055 33.165 165.065 ;
        RECT 34.475 155.055 34.745 165.065 ;
        RECT 36.055 155.055 36.325 165.065 ;
        RECT 106.745 155.055 107.015 165.065 ;
        RECT 108.325 155.055 108.595 165.065 ;
        RECT 109.905 155.055 110.175 165.065 ;
        RECT 111.485 155.055 111.755 165.065 ;
        RECT 113.065 155.055 113.335 165.065 ;
        RECT 114.645 155.055 114.915 165.065 ;
        RECT 116.225 155.055 116.495 165.065 ;
        RECT 117.805 155.055 118.075 165.065 ;
        RECT 119.385 155.055 119.655 165.065 ;
        RECT 34.585 154.165 35.765 154.215 ;
        RECT 107.305 154.165 108.485 154.215 ;
        RECT 120.835 154.165 121.125 165.955 ;
        RECT 21.945 153.935 37.795 154.165 ;
        RECT 105.275 153.935 121.125 154.165 ;
        RECT 34.585 153.885 35.765 153.935 ;
        RECT 107.305 153.885 108.485 153.935 ;
        RECT 23.265 146.535 23.535 151.535 ;
        RECT 24.845 146.535 25.115 151.535 ;
        RECT 26.425 146.535 26.695 151.535 ;
        RECT 28.005 146.535 28.275 151.535 ;
        RECT 29.585 146.535 29.855 151.535 ;
        RECT 31.165 146.535 31.435 151.535 ;
        RECT 35.025 150.625 35.255 151.285 ;
        RECT 36.605 150.625 36.835 151.285 ;
        RECT 35.025 149.745 36.835 150.625 ;
        RECT 35.025 149.085 35.255 149.745 ;
        RECT 36.605 149.085 36.835 149.745 ;
        RECT 106.235 150.625 106.465 151.285 ;
        RECT 107.815 150.625 108.045 151.285 ;
        RECT 106.235 149.745 108.045 150.625 ;
        RECT 106.235 149.085 106.465 149.745 ;
        RECT 107.815 149.085 108.045 149.745 ;
        RECT 111.635 146.535 111.905 151.535 ;
        RECT 113.215 146.535 113.485 151.535 ;
        RECT 114.795 146.535 115.065 151.535 ;
        RECT 116.375 146.535 116.645 151.535 ;
        RECT 117.955 146.535 118.225 151.535 ;
        RECT 119.535 146.535 119.805 151.535 ;
        RECT 20.750 144.945 21.910 144.965 ;
        RECT 19.590 144.915 21.910 144.945 ;
        RECT 121.160 144.945 122.320 144.965 ;
        RECT 121.160 144.915 123.480 144.945 ;
        RECT 19.590 143.995 22.240 144.915 ;
        RECT 120.830 143.995 123.480 144.915 ;
        RECT 19.590 143.965 21.910 143.995 ;
        RECT 121.160 143.965 123.480 143.995 ;
        RECT 19.590 143.945 21.100 143.965 ;
        RECT 121.970 143.945 123.480 143.965 ;
        RECT 23.060 137.580 23.290 138.240 ;
        RECT 24.640 137.580 24.870 138.240 ;
        RECT 23.060 136.700 24.870 137.580 ;
        RECT 23.060 136.040 23.290 136.700 ;
        RECT 24.640 136.040 24.870 136.700 ;
        RECT 118.200 137.580 118.430 138.240 ;
        RECT 119.780 137.580 120.010 138.240 ;
        RECT 118.200 136.700 120.010 137.580 ;
        RECT 118.200 136.040 118.430 136.700 ;
        RECT 119.780 136.040 120.010 136.700 ;
        RECT 24.130 133.390 25.310 133.440 ;
        RECT 117.760 133.390 118.940 133.440 ;
        RECT 22.100 133.160 37.950 133.390 ;
        RECT 24.130 133.110 25.310 133.160 ;
        RECT 37.660 121.370 37.950 133.160 ;
        RECT 22.100 121.140 37.950 121.370 ;
        RECT 105.120 133.160 120.970 133.390 ;
        RECT 105.120 121.370 105.410 133.160 ;
        RECT 117.760 133.110 118.940 133.160 ;
        RECT 105.120 121.140 120.970 121.370 ;
        RECT 22.605 117.725 38.455 117.955 ;
        RECT 22.605 105.935 22.895 117.725 ;
        RECT 105.275 117.055 121.125 117.285 ;
        RECT 24.075 106.825 24.345 116.835 ;
        RECT 25.655 106.825 25.925 116.835 ;
        RECT 27.235 106.825 27.505 116.835 ;
        RECT 28.815 106.825 29.085 116.835 ;
        RECT 30.395 106.825 30.665 116.835 ;
        RECT 31.975 106.825 32.245 116.835 ;
        RECT 33.555 106.825 33.825 116.835 ;
        RECT 35.135 106.825 35.405 116.835 ;
        RECT 36.715 106.825 36.985 116.835 ;
        RECT 106.745 106.155 107.015 116.165 ;
        RECT 108.325 106.155 108.595 116.165 ;
        RECT 109.905 106.155 110.175 116.165 ;
        RECT 111.485 106.155 111.755 116.165 ;
        RECT 113.065 106.155 113.335 116.165 ;
        RECT 114.645 106.155 114.915 116.165 ;
        RECT 116.225 106.155 116.495 116.165 ;
        RECT 117.805 106.155 118.075 116.165 ;
        RECT 119.385 106.155 119.655 116.165 ;
        RECT 35.245 105.935 36.425 105.985 ;
        RECT 22.605 105.705 38.455 105.935 ;
        RECT 35.245 105.655 36.425 105.705 ;
        RECT 107.305 105.265 108.485 105.315 ;
        RECT 120.835 105.265 121.125 117.055 ;
        RECT 105.275 105.035 121.125 105.265 ;
        RECT 107.305 104.985 108.485 105.035 ;
        RECT 23.925 98.305 24.195 103.305 ;
        RECT 25.505 98.305 25.775 103.305 ;
        RECT 27.085 98.305 27.355 103.305 ;
        RECT 28.665 98.305 28.935 103.305 ;
        RECT 30.245 98.305 30.515 103.305 ;
        RECT 31.825 98.305 32.095 103.305 ;
        RECT 35.685 102.395 35.915 103.055 ;
        RECT 37.265 102.395 37.495 103.055 ;
        RECT 35.685 101.515 37.495 102.395 ;
        RECT 35.685 100.855 35.915 101.515 ;
        RECT 37.265 100.855 37.495 101.515 ;
        RECT 106.235 101.725 106.465 102.385 ;
        RECT 107.815 101.725 108.045 102.385 ;
        RECT 106.235 100.845 108.045 101.725 ;
        RECT 106.235 100.185 106.465 100.845 ;
        RECT 107.815 100.185 108.045 100.845 ;
        RECT 111.635 97.635 111.905 102.635 ;
        RECT 113.215 97.635 113.485 102.635 ;
        RECT 114.795 97.635 115.065 102.635 ;
        RECT 116.375 97.635 116.645 102.635 ;
        RECT 117.955 97.635 118.225 102.635 ;
        RECT 119.535 97.635 119.805 102.635 ;
        RECT 21.410 96.715 22.570 96.735 ;
        RECT 20.250 96.685 22.570 96.715 ;
        RECT 20.250 95.765 22.900 96.685 ;
        RECT 121.160 96.045 122.320 96.065 ;
        RECT 121.160 96.015 123.480 96.045 ;
        RECT 20.250 95.735 22.570 95.765 ;
        RECT 20.250 95.715 21.760 95.735 ;
        RECT 120.830 95.095 123.480 96.015 ;
        RECT 121.160 95.065 123.480 95.095 ;
        RECT 121.970 95.045 123.480 95.065 ;
        RECT 23.720 89.350 23.950 90.010 ;
        RECT 25.300 89.350 25.530 90.010 ;
        RECT 23.720 88.470 25.530 89.350 ;
        RECT 23.720 87.810 23.950 88.470 ;
        RECT 25.300 87.810 25.530 88.470 ;
        RECT 118.200 88.680 118.430 89.340 ;
        RECT 119.780 88.680 120.010 89.340 ;
        RECT 118.200 87.800 120.010 88.680 ;
        RECT 118.200 87.140 118.430 87.800 ;
        RECT 119.780 87.140 120.010 87.800 ;
        RECT 24.790 85.160 25.970 85.210 ;
        RECT 22.760 84.930 38.610 85.160 ;
        RECT 24.790 84.880 25.970 84.930 ;
        RECT 38.320 73.140 38.610 84.930 ;
        RECT 117.760 84.490 118.940 84.540 ;
        RECT 22.760 72.910 38.610 73.140 ;
        RECT 105.120 84.260 120.970 84.490 ;
        RECT 105.120 72.470 105.410 84.260 ;
        RECT 117.760 84.210 118.940 84.260 ;
        RECT 105.120 72.240 120.970 72.470 ;
        RECT 22.275 67.155 38.125 67.385 ;
        RECT 104.615 67.155 120.465 67.385 ;
        RECT 22.275 55.365 22.565 67.155 ;
        RECT 23.745 56.255 24.015 66.265 ;
        RECT 25.325 56.255 25.595 66.265 ;
        RECT 26.905 56.255 27.175 66.265 ;
        RECT 28.485 56.255 28.755 66.265 ;
        RECT 30.065 56.255 30.335 66.265 ;
        RECT 31.645 56.255 31.915 66.265 ;
        RECT 33.225 56.255 33.495 66.265 ;
        RECT 34.805 56.255 35.075 66.265 ;
        RECT 36.385 56.255 36.655 66.265 ;
        RECT 106.085 56.255 106.355 66.265 ;
        RECT 107.665 56.255 107.935 66.265 ;
        RECT 109.245 56.255 109.515 66.265 ;
        RECT 110.825 56.255 111.095 66.265 ;
        RECT 112.405 56.255 112.675 66.265 ;
        RECT 113.985 56.255 114.255 66.265 ;
        RECT 115.565 56.255 115.835 66.265 ;
        RECT 117.145 56.255 117.415 66.265 ;
        RECT 118.725 56.255 118.995 66.265 ;
        RECT 34.915 55.365 36.095 55.415 ;
        RECT 106.645 55.365 107.825 55.415 ;
        RECT 120.175 55.365 120.465 67.155 ;
        RECT 22.275 55.135 38.125 55.365 ;
        RECT 104.615 55.135 120.465 55.365 ;
        RECT 34.915 55.085 36.095 55.135 ;
        RECT 106.645 55.085 107.825 55.135 ;
        RECT 23.595 47.735 23.865 52.735 ;
        RECT 25.175 47.735 25.445 52.735 ;
        RECT 26.755 47.735 27.025 52.735 ;
        RECT 28.335 47.735 28.605 52.735 ;
        RECT 29.915 47.735 30.185 52.735 ;
        RECT 31.495 47.735 31.765 52.735 ;
        RECT 35.355 51.825 35.585 52.485 ;
        RECT 36.935 51.825 37.165 52.485 ;
        RECT 35.355 50.945 37.165 51.825 ;
        RECT 35.355 50.285 35.585 50.945 ;
        RECT 36.935 50.285 37.165 50.945 ;
        RECT 105.575 51.825 105.805 52.485 ;
        RECT 107.155 51.825 107.385 52.485 ;
        RECT 105.575 50.945 107.385 51.825 ;
        RECT 105.575 50.285 105.805 50.945 ;
        RECT 107.155 50.285 107.385 50.945 ;
        RECT 110.975 47.735 111.245 52.735 ;
        RECT 112.555 47.735 112.825 52.735 ;
        RECT 114.135 47.735 114.405 52.735 ;
        RECT 115.715 47.735 115.985 52.735 ;
        RECT 117.295 47.735 117.565 52.735 ;
        RECT 118.875 47.735 119.145 52.735 ;
        RECT 21.080 46.145 22.240 46.165 ;
        RECT 19.920 46.115 22.240 46.145 ;
        RECT 120.500 46.145 121.660 46.165 ;
        RECT 120.500 46.115 122.820 46.145 ;
        RECT 19.920 45.195 22.570 46.115 ;
        RECT 120.170 45.195 122.820 46.115 ;
        RECT 19.920 45.165 22.240 45.195 ;
        RECT 120.500 45.165 122.820 45.195 ;
        RECT 19.920 45.145 21.430 45.165 ;
        RECT 121.310 45.145 122.820 45.165 ;
        RECT 23.390 38.780 23.620 39.440 ;
        RECT 24.970 38.780 25.200 39.440 ;
        RECT 23.390 37.900 25.200 38.780 ;
        RECT 23.390 37.240 23.620 37.900 ;
        RECT 24.970 37.240 25.200 37.900 ;
        RECT 117.540 38.780 117.770 39.440 ;
        RECT 119.120 38.780 119.350 39.440 ;
        RECT 117.540 37.900 119.350 38.780 ;
        RECT 117.540 37.240 117.770 37.900 ;
        RECT 119.120 37.240 119.350 37.900 ;
        RECT 24.460 34.590 25.640 34.640 ;
        RECT 117.100 34.590 118.280 34.640 ;
        RECT 22.430 34.360 38.280 34.590 ;
        RECT 24.460 34.310 25.640 34.360 ;
        RECT 37.990 22.570 38.280 34.360 ;
        RECT 22.430 22.340 38.280 22.570 ;
        RECT 104.460 34.360 120.310 34.590 ;
        RECT 104.460 22.570 104.750 34.360 ;
        RECT 117.100 34.310 118.280 34.360 ;
        RECT 104.460 22.340 120.310 22.570 ;
      LAYER met2 ;
        RECT 23.415 209.965 39.075 211.965 ;
        RECT 37.615 206.625 39.075 209.965 ;
        RECT 23.415 204.625 39.075 206.625 ;
        RECT 103.995 209.965 119.655 211.965 ;
        RECT 103.995 206.625 105.455 209.965 ;
        RECT 103.995 204.625 119.655 206.625 ;
        RECT 34.585 203.455 35.765 203.785 ;
        RECT 107.305 203.455 108.485 203.785 ;
        RECT 23.265 199.105 31.435 201.105 ;
        RECT 35.025 199.315 36.835 200.195 ;
        RECT 106.235 199.315 108.045 200.195 ;
        RECT 111.635 199.105 119.805 201.105 ;
        RECT 20.750 194.455 21.250 194.535 ;
        RECT 121.820 194.455 122.320 194.535 ;
        RECT 20.750 193.585 21.770 194.455 ;
        RECT 121.300 193.585 122.320 194.455 ;
        RECT 20.750 193.545 21.250 193.585 ;
        RECT 121.820 193.545 122.320 193.585 ;
        RECT 23.060 186.270 24.870 187.150 ;
        RECT 118.200 186.270 120.010 187.150 ;
        RECT 24.130 182.680 25.310 183.010 ;
        RECT 117.760 182.680 118.940 183.010 ;
        RECT 23.415 160.395 39.075 162.395 ;
        RECT 37.615 157.055 39.075 160.395 ;
        RECT 23.415 155.055 39.075 157.055 ;
        RECT 103.995 160.395 119.655 162.395 ;
        RECT 103.995 157.055 105.455 160.395 ;
        RECT 103.995 155.055 119.655 157.055 ;
        RECT 34.585 153.885 35.765 154.215 ;
        RECT 107.305 153.885 108.485 154.215 ;
        RECT 23.265 149.535 31.435 151.535 ;
        RECT 35.025 149.745 36.835 150.625 ;
        RECT 106.235 149.745 108.045 150.625 ;
        RECT 111.635 149.535 119.805 151.535 ;
        RECT 20.750 144.885 21.250 144.965 ;
        RECT 121.820 144.885 122.320 144.965 ;
        RECT 20.750 144.015 21.770 144.885 ;
        RECT 121.300 144.015 122.320 144.885 ;
        RECT 20.750 143.975 21.250 144.015 ;
        RECT 121.820 143.975 122.320 144.015 ;
        RECT 23.060 136.700 24.870 137.580 ;
        RECT 118.200 136.700 120.010 137.580 ;
        RECT 24.130 133.110 25.310 133.440 ;
        RECT 117.760 133.110 118.940 133.440 ;
        RECT 24.075 112.165 39.735 114.165 ;
        RECT 38.275 108.825 39.735 112.165 ;
        RECT 24.075 106.825 39.735 108.825 ;
        RECT 103.995 111.495 119.655 113.495 ;
        RECT 103.995 108.155 105.455 111.495 ;
        RECT 103.995 106.155 119.655 108.155 ;
        RECT 35.245 105.655 36.425 105.985 ;
        RECT 107.305 104.985 108.485 105.315 ;
        RECT 23.925 101.305 32.095 103.305 ;
        RECT 35.685 101.515 37.495 102.395 ;
        RECT 106.235 100.845 108.045 101.725 ;
        RECT 111.635 100.635 119.805 102.635 ;
        RECT 21.410 96.655 21.910 96.735 ;
        RECT 21.410 95.785 22.430 96.655 ;
        RECT 121.820 95.985 122.320 96.065 ;
        RECT 21.410 95.745 21.910 95.785 ;
        RECT 121.300 95.115 122.320 95.985 ;
        RECT 121.820 95.075 122.320 95.115 ;
        RECT 23.720 88.470 25.530 89.350 ;
        RECT 118.200 87.800 120.010 88.680 ;
        RECT 24.790 84.880 25.970 85.210 ;
        RECT 117.760 84.210 118.940 84.540 ;
        RECT 23.745 61.595 39.405 63.595 ;
        RECT 37.945 58.255 39.405 61.595 ;
        RECT 23.745 56.255 39.405 58.255 ;
        RECT 103.335 61.595 118.995 63.595 ;
        RECT 103.335 58.255 104.795 61.595 ;
        RECT 103.335 56.255 118.995 58.255 ;
        RECT 34.915 55.085 36.095 55.415 ;
        RECT 106.645 55.085 107.825 55.415 ;
        RECT 23.595 50.735 31.765 52.735 ;
        RECT 35.355 50.945 37.165 51.825 ;
        RECT 105.575 50.945 107.385 51.825 ;
        RECT 110.975 50.735 119.145 52.735 ;
        RECT 21.080 46.085 21.580 46.165 ;
        RECT 121.160 46.085 121.660 46.165 ;
        RECT 21.080 45.215 22.100 46.085 ;
        RECT 120.640 45.215 121.660 46.085 ;
        RECT 21.080 45.175 21.580 45.215 ;
        RECT 121.160 45.175 121.660 45.215 ;
        RECT 23.390 37.900 25.200 38.780 ;
        RECT 117.540 37.900 119.350 38.780 ;
        RECT 24.460 34.310 25.640 34.640 ;
        RECT 117.100 34.310 118.280 34.640 ;
      LAYER met3 ;
        RECT 23.415 204.625 39.075 206.625 ;
        RECT 103.995 204.625 119.655 206.625 ;
        RECT 28.875 203.095 30.875 204.625 ;
        RECT 34.585 203.425 35.765 203.815 ;
        RECT 107.305 203.425 108.485 203.815 ;
        RECT 112.195 203.095 114.195 204.625 ;
        RECT 28.875 202.435 34.490 203.095 ;
        RECT 108.580 202.435 114.195 203.095 ;
        RECT 28.875 201.105 30.875 202.435 ;
        RECT 24.015 199.105 31.435 201.105 ;
        RECT 33.240 195.855 34.230 202.435 ;
        RECT 34.575 199.315 36.835 200.195 ;
        RECT 106.235 199.315 108.495 200.195 ;
        RECT 108.840 195.855 109.830 202.435 ;
        RECT 112.195 201.105 114.195 202.435 ;
        RECT 111.635 199.105 119.055 201.105 ;
        RECT 33.240 195.355 34.020 195.855 ;
        RECT 109.050 195.355 109.830 195.855 ;
        RECT 20.610 194.575 21.950 194.635 ;
        RECT 20.610 194.495 23.170 194.575 ;
        RECT 33.240 194.495 33.970 195.355 ;
        RECT 109.100 194.495 109.830 195.355 ;
        RECT 121.120 194.575 122.460 194.635 ;
        RECT 119.900 194.495 122.460 194.575 ;
        RECT 20.610 194.475 33.970 194.495 ;
        RECT 20.610 194.325 34.020 194.475 ;
        RECT 20.610 194.295 34.060 194.325 ;
        RECT 20.610 194.285 34.240 194.295 ;
        RECT 34.950 194.285 35.740 194.495 ;
        RECT 20.610 193.455 35.740 194.285 ;
        RECT 21.830 193.395 35.740 193.455 ;
        RECT 107.330 194.285 108.120 194.495 ;
        RECT 109.100 194.475 122.460 194.495 ;
        RECT 109.050 194.325 122.460 194.475 ;
        RECT 109.010 194.295 122.460 194.325 ;
        RECT 108.830 194.285 122.460 194.295 ;
        RECT 107.330 193.455 122.460 194.285 ;
        RECT 107.330 193.395 121.240 193.455 ;
        RECT 23.060 186.270 25.320 187.150 ;
        RECT 117.750 186.270 120.010 187.150 ;
        RECT 24.130 182.650 25.310 183.040 ;
        RECT 117.760 182.650 118.940 183.040 ;
        RECT 23.415 155.055 39.075 157.055 ;
        RECT 103.995 155.055 119.655 157.055 ;
        RECT 28.875 153.525 30.875 155.055 ;
        RECT 34.585 153.855 35.765 154.245 ;
        RECT 107.305 153.855 108.485 154.245 ;
        RECT 112.195 153.525 114.195 155.055 ;
        RECT 28.875 152.865 34.490 153.525 ;
        RECT 108.580 152.865 114.195 153.525 ;
        RECT 28.875 151.535 30.875 152.865 ;
        RECT 24.015 149.535 31.435 151.535 ;
        RECT 33.240 146.285 34.230 152.865 ;
        RECT 34.575 149.745 36.835 150.625 ;
        RECT 106.235 149.745 108.495 150.625 ;
        RECT 108.840 146.285 109.830 152.865 ;
        RECT 112.195 151.535 114.195 152.865 ;
        RECT 111.635 149.535 119.055 151.535 ;
        RECT 33.240 145.785 34.020 146.285 ;
        RECT 109.050 145.785 109.830 146.285 ;
        RECT 20.610 145.005 21.950 145.065 ;
        RECT 20.610 144.925 23.170 145.005 ;
        RECT 33.240 144.925 33.970 145.785 ;
        RECT 109.100 144.925 109.830 145.785 ;
        RECT 121.120 145.005 122.460 145.065 ;
        RECT 119.900 144.925 122.460 145.005 ;
        RECT 20.610 144.905 33.970 144.925 ;
        RECT 20.610 144.755 34.020 144.905 ;
        RECT 20.610 144.725 34.060 144.755 ;
        RECT 20.610 144.715 34.240 144.725 ;
        RECT 34.950 144.715 35.740 144.925 ;
        RECT 20.610 143.885 35.740 144.715 ;
        RECT 21.830 143.825 35.740 143.885 ;
        RECT 107.330 144.715 108.120 144.925 ;
        RECT 109.100 144.905 122.460 144.925 ;
        RECT 109.050 144.755 122.460 144.905 ;
        RECT 109.010 144.725 122.460 144.755 ;
        RECT 108.830 144.715 122.460 144.725 ;
        RECT 107.330 143.885 122.460 144.715 ;
        RECT 107.330 143.825 121.240 143.885 ;
        RECT 23.060 136.700 25.320 137.580 ;
        RECT 117.750 136.700 120.010 137.580 ;
        RECT 24.130 133.080 25.310 133.470 ;
        RECT 117.760 133.080 118.940 133.470 ;
        RECT 24.075 106.825 39.735 108.825 ;
        RECT 29.535 105.295 31.535 106.825 ;
        RECT 103.995 106.155 119.655 108.155 ;
        RECT 35.245 105.625 36.425 106.015 ;
        RECT 29.535 104.635 35.150 105.295 ;
        RECT 107.305 104.955 108.485 105.345 ;
        RECT 29.535 103.305 31.535 104.635 ;
        RECT 24.675 101.305 32.095 103.305 ;
        RECT 33.900 98.055 34.890 104.635 ;
        RECT 112.195 104.625 114.195 106.155 ;
        RECT 108.580 103.965 114.195 104.625 ;
        RECT 35.235 101.515 37.495 102.395 ;
        RECT 106.235 100.845 108.495 101.725 ;
        RECT 33.900 97.555 34.680 98.055 ;
        RECT 21.270 96.775 22.610 96.835 ;
        RECT 21.270 96.695 23.830 96.775 ;
        RECT 33.900 96.695 34.630 97.555 ;
        RECT 108.840 97.385 109.830 103.965 ;
        RECT 112.195 102.635 114.195 103.965 ;
        RECT 111.635 100.635 119.055 102.635 ;
        RECT 109.050 96.885 109.830 97.385 ;
        RECT 21.270 96.675 34.630 96.695 ;
        RECT 21.270 96.525 34.680 96.675 ;
        RECT 21.270 96.495 34.720 96.525 ;
        RECT 21.270 96.485 34.900 96.495 ;
        RECT 35.610 96.485 36.400 96.695 ;
        RECT 21.270 95.655 36.400 96.485 ;
        RECT 109.100 96.025 109.830 96.885 ;
        RECT 121.120 96.105 122.460 96.165 ;
        RECT 119.900 96.025 122.460 96.105 ;
        RECT 22.490 95.595 36.400 95.655 ;
        RECT 107.330 95.815 108.120 96.025 ;
        RECT 109.100 96.005 122.460 96.025 ;
        RECT 109.050 95.855 122.460 96.005 ;
        RECT 109.010 95.825 122.460 95.855 ;
        RECT 108.830 95.815 122.460 95.825 ;
        RECT 107.330 94.985 122.460 95.815 ;
        RECT 107.330 94.925 121.240 94.985 ;
        RECT 23.720 88.470 25.980 89.350 ;
        RECT 117.750 87.800 120.010 88.680 ;
        RECT 24.790 84.850 25.970 85.240 ;
        RECT 117.760 84.180 118.940 84.570 ;
        RECT 23.745 56.255 39.405 58.255 ;
        RECT 103.335 56.255 118.995 58.255 ;
        RECT 29.205 54.725 31.205 56.255 ;
        RECT 34.915 55.055 36.095 55.445 ;
        RECT 106.645 55.055 107.825 55.445 ;
        RECT 111.535 54.725 113.535 56.255 ;
        RECT 29.205 54.065 34.820 54.725 ;
        RECT 107.920 54.065 113.535 54.725 ;
        RECT 29.205 52.735 31.205 54.065 ;
        RECT 24.345 50.735 31.765 52.735 ;
        RECT 33.570 47.485 34.560 54.065 ;
        RECT 34.905 50.945 37.165 51.825 ;
        RECT 105.575 50.945 107.835 51.825 ;
        RECT 108.180 47.485 109.170 54.065 ;
        RECT 111.535 52.735 113.535 54.065 ;
        RECT 110.975 50.735 118.395 52.735 ;
        RECT 33.570 46.985 34.350 47.485 ;
        RECT 108.390 46.985 109.170 47.485 ;
        RECT 20.940 46.205 22.280 46.265 ;
        RECT 20.940 46.125 23.500 46.205 ;
        RECT 33.570 46.125 34.300 46.985 ;
        RECT 108.440 46.125 109.170 46.985 ;
        RECT 120.460 46.205 121.800 46.265 ;
        RECT 119.240 46.125 121.800 46.205 ;
        RECT 20.940 46.105 34.300 46.125 ;
        RECT 20.940 45.955 34.350 46.105 ;
        RECT 20.940 45.925 34.390 45.955 ;
        RECT 20.940 45.915 34.570 45.925 ;
        RECT 35.280 45.915 36.070 46.125 ;
        RECT 20.940 45.085 36.070 45.915 ;
        RECT 22.160 45.025 36.070 45.085 ;
        RECT 106.670 45.915 107.460 46.125 ;
        RECT 108.440 46.105 121.800 46.125 ;
        RECT 108.390 45.955 121.800 46.105 ;
        RECT 108.350 45.925 121.800 45.955 ;
        RECT 108.170 45.915 121.800 45.925 ;
        RECT 106.670 45.085 121.800 45.915 ;
        RECT 106.670 45.025 120.580 45.085 ;
        RECT 23.390 37.900 25.650 38.780 ;
        RECT 117.090 37.900 119.350 38.780 ;
        RECT 24.460 34.280 25.640 34.670 ;
        RECT 117.100 34.280 118.280 34.670 ;
      LAYER met4 ;
        RECT 7.000 194.400 9.000 220.760 ;
        RECT 29.425 202.605 30.325 204.605 ;
        RECT 34.575 194.675 35.775 216.365 ;
        RECT 34.550 194.605 35.775 194.675 ;
        RECT 107.295 194.675 108.495 216.365 ;
        RECT 112.745 202.605 113.645 204.605 ;
        RECT 107.295 194.605 108.520 194.675 ;
        RECT 7.000 194.375 18.660 194.400 ;
        RECT 24.060 194.375 25.250 194.495 ;
        RECT 7.000 193.570 25.290 194.375 ;
        RECT 7.000 144.850 9.000 193.570 ;
        RECT 18.040 193.535 25.290 193.570 ;
        RECT 24.060 191.860 25.250 193.535 ;
        RECT 34.550 193.375 35.730 194.605 ;
        RECT 107.340 193.375 108.520 194.605 ;
        RECT 117.820 194.375 119.010 194.495 ;
        RECT 131.865 194.375 133.920 223.215 ;
        RECT 117.780 193.535 133.920 194.375 ;
        RECT 117.820 191.860 119.010 193.535 ;
        RECT 24.060 191.705 25.320 191.860 ;
        RECT 24.120 170.100 25.320 191.705 ;
        RECT 117.750 191.705 119.010 191.860 ;
        RECT 117.750 170.100 118.950 191.705 ;
        RECT 29.425 153.035 30.325 155.035 ;
        RECT 34.575 145.105 35.775 166.795 ;
        RECT 34.550 145.035 35.775 145.105 ;
        RECT 107.295 145.105 108.495 166.795 ;
        RECT 112.745 153.035 113.645 155.035 ;
        RECT 107.295 145.035 108.520 145.105 ;
        RECT 7.000 144.805 18.850 144.850 ;
        RECT 24.060 144.805 25.250 144.925 ;
        RECT 7.000 143.990 25.290 144.805 ;
        RECT 7.000 115.400 9.000 143.990 ;
        RECT 18.040 143.965 25.290 143.990 ;
        RECT 24.060 142.290 25.250 143.965 ;
        RECT 34.550 143.805 35.730 145.035 ;
        RECT 107.340 143.805 108.520 145.035 ;
        RECT 117.820 144.805 119.010 144.925 ;
        RECT 131.865 144.805 133.920 193.535 ;
        RECT 117.780 143.965 133.920 144.805 ;
        RECT 117.820 142.290 119.010 143.965 ;
        RECT 24.060 142.135 25.320 142.290 ;
        RECT 24.120 120.530 25.320 142.135 ;
        RECT 117.750 142.135 119.010 142.290 ;
        RECT 117.750 120.530 118.950 142.135 ;
        RECT 7.000 112.600 9.030 115.400 ;
        RECT 7.000 103.450 9.000 112.600 ;
        RECT 30.085 104.805 30.985 106.805 ;
        RECT 7.000 101.970 9.050 103.450 ;
        RECT 7.000 96.510 9.000 101.970 ;
        RECT 35.235 96.875 36.435 118.565 ;
        RECT 35.210 96.805 36.435 96.875 ;
        RECT 24.720 96.575 25.910 96.695 ;
        RECT 18.700 96.510 25.950 96.575 ;
        RECT 6.980 95.735 25.950 96.510 ;
        RECT 6.980 95.650 18.830 95.735 ;
        RECT 7.000 69.170 9.000 95.650 ;
        RECT 24.720 94.060 25.910 95.735 ;
        RECT 35.210 95.575 36.390 96.805 ;
        RECT 107.295 96.205 108.495 117.895 ;
        RECT 112.745 104.135 113.645 106.135 ;
        RECT 107.295 96.135 108.520 96.205 ;
        RECT 107.340 94.905 108.520 96.135 ;
        RECT 117.820 95.905 119.010 96.025 ;
        RECT 131.865 95.905 133.920 143.965 ;
        RECT 117.780 95.065 133.920 95.905 ;
        RECT 24.720 93.905 25.980 94.060 ;
        RECT 24.780 72.300 25.980 93.905 ;
        RECT 117.820 93.390 119.010 95.065 ;
        RECT 117.750 93.235 119.010 93.390 ;
        RECT 117.750 71.630 118.950 93.235 ;
        RECT 7.000 67.690 9.010 69.170 ;
        RECT 7.000 46.040 9.000 67.690 ;
        RECT 29.755 54.235 30.655 56.235 ;
        RECT 34.905 46.305 36.105 67.995 ;
        RECT 34.880 46.235 36.105 46.305 ;
        RECT 106.635 46.305 107.835 67.995 ;
        RECT 112.085 54.235 112.985 56.235 ;
        RECT 106.635 46.235 107.860 46.305 ;
        RECT 7.000 46.005 18.880 46.040 ;
        RECT 24.390 46.005 25.580 46.125 ;
        RECT 7.000 45.180 25.620 46.005 ;
        RECT 7.000 13.950 9.000 45.180 ;
        RECT 18.370 45.165 25.620 45.180 ;
        RECT 24.390 43.490 25.580 45.165 ;
        RECT 34.880 45.005 36.060 46.235 ;
        RECT 106.680 45.005 107.860 46.235 ;
        RECT 117.160 46.005 118.350 46.125 ;
        RECT 131.865 46.005 133.920 95.065 ;
        RECT 117.120 45.165 133.920 46.005 ;
        RECT 117.160 43.490 118.350 45.165 ;
        RECT 24.390 43.335 25.650 43.490 ;
        RECT 24.450 21.730 25.650 43.335 ;
        RECT 117.090 43.335 118.350 43.490 ;
        RECT 41.490 26.640 46.490 27.790 ;
        RECT 41.110 17.790 46.490 26.640 ;
        RECT 117.090 21.730 118.290 43.335 ;
        RECT 41.110 13.950 46.290 17.790 ;
        RECT 131.865 13.950 133.920 45.165 ;
        RECT 7.000 11.940 133.920 13.950 ;
        RECT 7.000 5.000 9.000 11.940 ;
        RECT 41.110 11.330 46.290 11.940 ;
        RECT 131.865 11.920 133.920 11.940 ;
    END
  END VAPWR
  OBS
      LAYER pwell ;
        RECT 15.515 186.785 16.425 187.820 ;
        RECT 15.325 186.615 16.425 186.785 ;
        RECT 15.515 186.470 16.425 186.615 ;
        RECT 126.645 186.785 127.555 187.820 ;
        RECT 126.645 186.615 127.745 186.785 ;
        RECT 126.645 186.470 127.555 186.615 ;
        RECT 15.250 183.110 16.180 184.020 ;
        RECT 16.970 183.110 17.900 184.020 ;
        RECT 16.075 183.090 16.180 183.110 ;
        RECT 17.795 183.090 17.900 183.110 ;
        RECT 125.170 183.110 126.100 184.020 ;
        RECT 126.890 183.110 127.820 184.020 ;
        RECT 125.170 183.090 125.275 183.110 ;
        RECT 126.890 183.090 126.995 183.110 ;
        RECT 16.075 182.920 16.245 183.090 ;
        RECT 17.795 182.920 17.965 183.090 ;
        RECT 125.105 182.920 125.275 183.090 ;
        RECT 126.825 182.920 126.995 183.090 ;
        RECT 15.410 179.000 16.340 179.910 ;
        RECT 17.070 179.010 18.000 179.920 ;
        RECT 16.235 178.980 16.340 179.000 ;
        RECT 17.895 178.990 18.000 179.010 ;
        RECT 125.070 179.010 126.000 179.920 ;
        RECT 125.070 178.990 125.175 179.010 ;
        RECT 16.235 178.810 16.405 178.980 ;
        RECT 17.895 178.820 18.065 178.990 ;
        RECT 125.005 178.820 125.175 178.990 ;
        RECT 126.730 179.000 127.660 179.910 ;
        RECT 126.730 178.980 126.835 179.000 ;
        RECT 126.665 178.810 126.835 178.980 ;
        RECT 15.445 177.015 16.355 178.050 ;
        RECT 15.255 176.845 16.355 177.015 ;
        RECT 15.445 176.700 16.355 176.845 ;
        RECT 126.715 177.015 127.625 178.050 ;
        RECT 126.715 176.845 127.815 177.015 ;
        RECT 126.715 176.700 127.625 176.845 ;
        RECT 15.415 175.410 16.325 176.235 ;
        RECT 15.225 175.305 16.325 175.410 ;
        RECT 126.745 175.410 127.655 176.235 ;
        RECT 126.745 175.305 127.845 175.410 ;
        RECT 15.225 175.240 15.395 175.305 ;
        RECT 127.675 175.240 127.845 175.305 ;
        RECT 15.515 137.215 16.425 138.250 ;
        RECT 15.325 137.045 16.425 137.215 ;
        RECT 15.515 136.900 16.425 137.045 ;
        RECT 126.645 137.215 127.555 138.250 ;
        RECT 126.645 137.045 127.745 137.215 ;
        RECT 126.645 136.900 127.555 137.045 ;
        RECT 15.250 133.540 16.180 134.450 ;
        RECT 16.970 133.540 17.900 134.450 ;
        RECT 16.075 133.520 16.180 133.540 ;
        RECT 17.795 133.520 17.900 133.540 ;
        RECT 125.170 133.540 126.100 134.450 ;
        RECT 126.890 133.540 127.820 134.450 ;
        RECT 125.170 133.520 125.275 133.540 ;
        RECT 126.890 133.520 126.995 133.540 ;
        RECT 16.075 133.350 16.245 133.520 ;
        RECT 17.795 133.350 17.965 133.520 ;
        RECT 125.105 133.350 125.275 133.520 ;
        RECT 126.825 133.350 126.995 133.520 ;
        RECT 15.410 129.430 16.340 130.340 ;
        RECT 17.070 129.440 18.000 130.350 ;
        RECT 16.235 129.410 16.340 129.430 ;
        RECT 17.895 129.420 18.000 129.440 ;
        RECT 125.070 129.440 126.000 130.350 ;
        RECT 125.070 129.420 125.175 129.440 ;
        RECT 16.235 129.240 16.405 129.410 ;
        RECT 17.895 129.250 18.065 129.420 ;
        RECT 125.005 129.250 125.175 129.420 ;
        RECT 126.730 129.430 127.660 130.340 ;
        RECT 126.730 129.410 126.835 129.430 ;
        RECT 126.665 129.240 126.835 129.410 ;
        RECT 15.445 127.445 16.355 128.480 ;
        RECT 15.255 127.275 16.355 127.445 ;
        RECT 15.445 127.130 16.355 127.275 ;
        RECT 126.715 127.445 127.625 128.480 ;
        RECT 126.715 127.275 127.815 127.445 ;
        RECT 126.715 127.130 127.625 127.275 ;
        RECT 15.415 125.840 16.325 126.665 ;
        RECT 15.225 125.735 16.325 125.840 ;
        RECT 126.745 125.840 127.655 126.665 ;
        RECT 126.745 125.735 127.845 125.840 ;
        RECT 15.225 125.670 15.395 125.735 ;
        RECT 127.675 125.670 127.845 125.735 ;
        RECT 16.175 88.985 17.085 90.020 ;
        RECT 15.985 88.815 17.085 88.985 ;
        RECT 16.175 88.670 17.085 88.815 ;
        RECT 126.645 88.315 127.555 89.350 ;
        RECT 126.645 88.145 127.745 88.315 ;
        RECT 126.645 88.000 127.555 88.145 ;
        RECT 15.910 85.310 16.840 86.220 ;
        RECT 17.630 85.310 18.560 86.220 ;
        RECT 16.735 85.290 16.840 85.310 ;
        RECT 18.455 85.290 18.560 85.310 ;
        RECT 16.735 85.120 16.905 85.290 ;
        RECT 18.455 85.120 18.625 85.290 ;
        RECT 125.170 84.640 126.100 85.550 ;
        RECT 126.890 84.640 127.820 85.550 ;
        RECT 125.170 84.620 125.275 84.640 ;
        RECT 126.890 84.620 126.995 84.640 ;
        RECT 125.105 84.450 125.275 84.620 ;
        RECT 126.825 84.450 126.995 84.620 ;
        RECT 16.070 81.200 17.000 82.110 ;
        RECT 17.730 81.210 18.660 82.120 ;
        RECT 16.895 81.180 17.000 81.200 ;
        RECT 18.555 81.190 18.660 81.210 ;
        RECT 16.895 81.010 17.065 81.180 ;
        RECT 18.555 81.020 18.725 81.190 ;
        RECT 125.070 80.540 126.000 81.450 ;
        RECT 125.070 80.520 125.175 80.540 ;
        RECT 125.005 80.350 125.175 80.520 ;
        RECT 126.730 80.530 127.660 81.440 ;
        RECT 126.730 80.510 126.835 80.530 ;
        RECT 126.665 80.340 126.835 80.510 ;
        RECT 16.105 79.215 17.015 80.250 ;
        RECT 15.915 79.045 17.015 79.215 ;
        RECT 16.105 78.900 17.015 79.045 ;
        RECT 126.715 78.545 127.625 79.580 ;
        RECT 16.075 77.610 16.985 78.435 ;
        RECT 126.715 78.375 127.815 78.545 ;
        RECT 126.715 78.230 127.625 78.375 ;
        RECT 15.885 77.505 16.985 77.610 ;
        RECT 15.885 77.440 16.055 77.505 ;
        RECT 126.745 76.940 127.655 77.765 ;
        RECT 126.745 76.835 127.845 76.940 ;
        RECT 127.675 76.770 127.845 76.835 ;
        RECT 15.845 38.415 16.755 39.450 ;
        RECT 15.655 38.245 16.755 38.415 ;
        RECT 15.845 38.100 16.755 38.245 ;
        RECT 125.985 38.415 126.895 39.450 ;
        RECT 125.985 38.245 127.085 38.415 ;
        RECT 125.985 38.100 126.895 38.245 ;
        RECT 15.580 34.740 16.510 35.650 ;
        RECT 17.300 34.740 18.230 35.650 ;
        RECT 16.405 34.720 16.510 34.740 ;
        RECT 18.125 34.720 18.230 34.740 ;
        RECT 124.510 34.740 125.440 35.650 ;
        RECT 126.230 34.740 127.160 35.650 ;
        RECT 124.510 34.720 124.615 34.740 ;
        RECT 126.230 34.720 126.335 34.740 ;
        RECT 16.405 34.550 16.575 34.720 ;
        RECT 18.125 34.550 18.295 34.720 ;
        RECT 124.445 34.550 124.615 34.720 ;
        RECT 126.165 34.550 126.335 34.720 ;
        RECT 15.740 30.630 16.670 31.540 ;
        RECT 17.400 30.640 18.330 31.550 ;
        RECT 16.565 30.610 16.670 30.630 ;
        RECT 18.225 30.620 18.330 30.640 ;
        RECT 124.410 30.640 125.340 31.550 ;
        RECT 124.410 30.620 124.515 30.640 ;
        RECT 16.565 30.440 16.735 30.610 ;
        RECT 18.225 30.450 18.395 30.620 ;
        RECT 124.345 30.450 124.515 30.620 ;
        RECT 126.070 30.630 127.000 31.540 ;
        RECT 126.070 30.610 126.175 30.630 ;
        RECT 126.005 30.440 126.175 30.610 ;
        RECT 15.775 28.645 16.685 29.680 ;
        RECT 15.585 28.475 16.685 28.645 ;
        RECT 15.775 28.330 16.685 28.475 ;
        RECT 126.055 28.645 126.965 29.680 ;
        RECT 126.055 28.475 127.155 28.645 ;
        RECT 126.055 28.330 126.965 28.475 ;
        RECT 15.745 27.040 16.655 27.865 ;
        RECT 15.555 26.935 16.655 27.040 ;
        RECT 126.085 27.040 126.995 27.865 ;
        RECT 126.085 26.935 127.185 27.040 ;
        RECT 15.555 26.870 15.725 26.935 ;
        RECT 127.015 26.870 127.185 26.935 ;
      LAYER li1 ;
        RECT 22.905 214.865 23.405 215.035 ;
        RECT 23.695 214.865 24.195 215.035 ;
        RECT 24.485 214.865 24.985 215.035 ;
        RECT 25.275 214.865 25.775 215.035 ;
        RECT 26.065 214.865 26.565 215.035 ;
        RECT 26.855 214.865 27.355 215.035 ;
        RECT 27.645 214.865 28.145 215.035 ;
        RECT 28.435 214.865 28.935 215.035 ;
        RECT 29.225 214.865 29.725 215.035 ;
        RECT 30.015 214.865 30.515 215.035 ;
        RECT 30.805 214.865 31.305 215.035 ;
        RECT 31.595 214.865 32.095 215.035 ;
        RECT 32.385 214.865 32.885 215.035 ;
        RECT 33.175 214.865 33.675 215.035 ;
        RECT 33.965 214.865 34.465 215.035 ;
        RECT 34.755 214.865 35.255 215.035 ;
        RECT 35.545 214.865 36.045 215.035 ;
        RECT 36.335 214.865 36.835 215.035 ;
        RECT 106.235 214.865 106.735 215.035 ;
        RECT 107.025 214.865 107.525 215.035 ;
        RECT 107.815 214.865 108.315 215.035 ;
        RECT 108.605 214.865 109.105 215.035 ;
        RECT 109.395 214.865 109.895 215.035 ;
        RECT 110.185 214.865 110.685 215.035 ;
        RECT 110.975 214.865 111.475 215.035 ;
        RECT 111.765 214.865 112.265 215.035 ;
        RECT 112.555 214.865 113.055 215.035 ;
        RECT 113.345 214.865 113.845 215.035 ;
        RECT 114.135 214.865 114.635 215.035 ;
        RECT 114.925 214.865 115.425 215.035 ;
        RECT 115.715 214.865 116.215 215.035 ;
        RECT 116.505 214.865 117.005 215.035 ;
        RECT 117.295 214.865 117.795 215.035 ;
        RECT 118.085 214.865 118.585 215.035 ;
        RECT 118.875 214.865 119.375 215.035 ;
        RECT 119.665 214.865 120.165 215.035 ;
        RECT 22.675 204.610 22.845 214.650 ;
        RECT 24.255 204.610 24.425 214.650 ;
        RECT 25.835 204.610 26.005 214.650 ;
        RECT 27.415 204.610 27.585 214.650 ;
        RECT 28.995 204.610 29.165 214.650 ;
        RECT 30.575 204.610 30.745 214.650 ;
        RECT 32.155 204.610 32.325 214.650 ;
        RECT 33.735 204.610 33.905 214.650 ;
        RECT 35.315 204.610 35.485 214.650 ;
        RECT 36.895 204.610 37.065 214.650 ;
        RECT 106.005 204.610 106.175 214.650 ;
        RECT 107.585 204.610 107.755 214.650 ;
        RECT 109.165 204.610 109.335 214.650 ;
        RECT 110.745 204.610 110.915 214.650 ;
        RECT 112.325 204.610 112.495 214.650 ;
        RECT 113.905 204.610 114.075 214.650 ;
        RECT 115.485 204.610 115.655 214.650 ;
        RECT 117.065 204.610 117.235 214.650 ;
        RECT 118.645 204.610 118.815 214.650 ;
        RECT 120.225 204.610 120.395 214.650 ;
        RECT 22.905 204.225 23.405 204.395 ;
        RECT 23.695 204.225 24.195 204.395 ;
        RECT 24.485 204.225 24.985 204.395 ;
        RECT 25.275 204.225 25.775 204.395 ;
        RECT 26.065 204.225 26.565 204.395 ;
        RECT 26.855 204.225 27.355 204.395 ;
        RECT 27.645 204.225 28.145 204.395 ;
        RECT 28.435 204.225 28.935 204.395 ;
        RECT 29.225 204.225 29.725 204.395 ;
        RECT 30.015 204.225 30.515 204.395 ;
        RECT 30.805 204.225 31.305 204.395 ;
        RECT 31.595 204.225 32.095 204.395 ;
        RECT 32.385 204.225 32.885 204.395 ;
        RECT 33.175 204.225 33.675 204.395 ;
        RECT 33.965 204.225 34.465 204.395 ;
        RECT 34.755 204.225 35.255 204.395 ;
        RECT 35.545 204.225 36.045 204.395 ;
        RECT 36.335 204.225 36.835 204.395 ;
        RECT 106.235 204.225 106.735 204.395 ;
        RECT 107.025 204.225 107.525 204.395 ;
        RECT 107.815 204.225 108.315 204.395 ;
        RECT 108.605 204.225 109.105 204.395 ;
        RECT 109.395 204.225 109.895 204.395 ;
        RECT 110.185 204.225 110.685 204.395 ;
        RECT 110.975 204.225 111.475 204.395 ;
        RECT 111.765 204.225 112.265 204.395 ;
        RECT 112.555 204.225 113.055 204.395 ;
        RECT 113.345 204.225 113.845 204.395 ;
        RECT 114.135 204.225 114.635 204.395 ;
        RECT 114.925 204.225 115.425 204.395 ;
        RECT 115.715 204.225 116.215 204.395 ;
        RECT 116.505 204.225 117.005 204.395 ;
        RECT 117.295 204.225 117.795 204.395 ;
        RECT 118.085 204.225 118.585 204.395 ;
        RECT 118.875 204.225 119.375 204.395 ;
        RECT 119.665 204.225 120.165 204.395 ;
        RECT 37.545 202.095 38.135 202.265 ;
        RECT 104.935 202.095 105.525 202.265 ;
        RECT 22.755 201.295 23.255 201.465 ;
        RECT 23.545 201.295 24.045 201.465 ;
        RECT 24.335 201.295 24.835 201.465 ;
        RECT 25.125 201.295 25.625 201.465 ;
        RECT 25.915 201.295 26.415 201.465 ;
        RECT 26.705 201.295 27.205 201.465 ;
        RECT 27.495 201.295 27.995 201.465 ;
        RECT 28.285 201.295 28.785 201.465 ;
        RECT 29.075 201.295 29.575 201.465 ;
        RECT 29.865 201.295 30.365 201.465 ;
        RECT 30.655 201.295 31.155 201.465 ;
        RECT 31.445 201.295 31.945 201.465 ;
        RECT 22.525 196.085 22.695 201.125 ;
        RECT 24.105 196.085 24.275 201.125 ;
        RECT 25.685 196.085 25.855 201.125 ;
        RECT 27.265 196.085 27.435 201.125 ;
        RECT 28.845 196.085 29.015 201.125 ;
        RECT 30.425 196.085 30.595 201.125 ;
        RECT 32.005 196.085 32.175 201.125 ;
        RECT 35.845 200.355 36.015 201.945 ;
        RECT 38.055 201.275 38.385 201.865 ;
        RECT 36.185 201.025 38.385 201.275 ;
        RECT 38.055 200.435 38.385 201.025 ;
        RECT 104.685 201.275 105.015 201.865 ;
        RECT 104.685 201.025 106.885 201.275 ;
        RECT 104.685 200.435 105.015 201.025 ;
        RECT 107.055 200.355 107.225 201.945 ;
        RECT 111.125 201.295 111.625 201.465 ;
        RECT 111.915 201.295 112.415 201.465 ;
        RECT 112.705 201.295 113.205 201.465 ;
        RECT 113.495 201.295 113.995 201.465 ;
        RECT 114.285 201.295 114.785 201.465 ;
        RECT 115.075 201.295 115.575 201.465 ;
        RECT 115.865 201.295 116.365 201.465 ;
        RECT 116.655 201.295 117.155 201.465 ;
        RECT 117.445 201.295 117.945 201.465 ;
        RECT 118.235 201.295 118.735 201.465 ;
        RECT 119.025 201.295 119.525 201.465 ;
        RECT 119.815 201.295 120.315 201.465 ;
        RECT 37.495 199.985 38.105 200.155 ;
        RECT 104.965 199.985 105.575 200.155 ;
        RECT 37.545 199.355 38.155 199.525 ;
        RECT 104.915 199.355 105.525 199.525 ;
        RECT 35.845 197.565 36.015 199.155 ;
        RECT 38.055 198.485 38.385 199.075 ;
        RECT 36.185 198.235 38.385 198.485 ;
        RECT 38.055 197.645 38.385 198.235 ;
        RECT 104.685 198.485 105.015 199.075 ;
        RECT 104.685 198.235 106.885 198.485 ;
        RECT 104.685 197.645 105.015 198.235 ;
        RECT 107.055 197.565 107.225 199.155 ;
        RECT 37.545 197.245 38.135 197.415 ;
        RECT 104.935 197.245 105.525 197.415 ;
        RECT 36.685 195.975 37.025 196.145 ;
        RECT 37.745 195.975 38.665 196.145 ;
        RECT 104.405 195.975 105.325 196.145 ;
        RECT 106.045 195.975 106.385 196.145 ;
        RECT 110.895 196.085 111.065 201.125 ;
        RECT 112.475 196.085 112.645 201.125 ;
        RECT 114.055 196.085 114.225 201.125 ;
        RECT 115.635 196.085 115.805 201.125 ;
        RECT 117.215 196.085 117.385 201.125 ;
        RECT 118.795 196.085 118.965 201.125 ;
        RECT 120.375 196.085 120.545 201.125 ;
        RECT 22.755 195.745 23.255 195.915 ;
        RECT 23.545 195.745 24.045 195.915 ;
        RECT 24.335 195.745 24.835 195.915 ;
        RECT 25.125 195.745 25.625 195.915 ;
        RECT 25.915 195.745 26.415 195.915 ;
        RECT 26.705 195.745 27.205 195.915 ;
        RECT 27.495 195.745 27.995 195.915 ;
        RECT 28.285 195.745 28.785 195.915 ;
        RECT 29.075 195.745 29.575 195.915 ;
        RECT 29.865 195.745 30.365 195.915 ;
        RECT 30.655 195.745 31.155 195.915 ;
        RECT 31.445 195.745 31.945 195.915 ;
        RECT 37.295 195.545 37.465 195.915 ;
        RECT 105.605 195.545 105.775 195.915 ;
        RECT 111.125 195.745 111.625 195.915 ;
        RECT 111.915 195.745 112.415 195.915 ;
        RECT 112.705 195.745 113.205 195.915 ;
        RECT 113.495 195.745 113.995 195.915 ;
        RECT 114.285 195.745 114.785 195.915 ;
        RECT 115.075 195.745 115.575 195.915 ;
        RECT 115.865 195.745 116.365 195.915 ;
        RECT 116.655 195.745 117.155 195.915 ;
        RECT 117.445 195.745 117.945 195.915 ;
        RECT 118.235 195.745 118.735 195.915 ;
        RECT 119.025 195.745 119.525 195.915 ;
        RECT 119.815 195.745 120.315 195.915 ;
        RECT 22.430 190.550 22.600 190.920 ;
        RECT 27.950 190.550 28.450 190.720 ;
        RECT 28.740 190.550 29.240 190.720 ;
        RECT 29.530 190.550 30.030 190.720 ;
        RECT 30.320 190.550 30.820 190.720 ;
        RECT 31.110 190.550 31.610 190.720 ;
        RECT 31.900 190.550 32.400 190.720 ;
        RECT 32.690 190.550 33.190 190.720 ;
        RECT 33.480 190.550 33.980 190.720 ;
        RECT 34.270 190.550 34.770 190.720 ;
        RECT 35.060 190.550 35.560 190.720 ;
        RECT 35.850 190.550 36.350 190.720 ;
        RECT 36.640 190.550 37.140 190.720 ;
        RECT 105.930 190.550 106.430 190.720 ;
        RECT 106.720 190.550 107.220 190.720 ;
        RECT 107.510 190.550 108.010 190.720 ;
        RECT 108.300 190.550 108.800 190.720 ;
        RECT 109.090 190.550 109.590 190.720 ;
        RECT 109.880 190.550 110.380 190.720 ;
        RECT 110.670 190.550 111.170 190.720 ;
        RECT 111.460 190.550 111.960 190.720 ;
        RECT 112.250 190.550 112.750 190.720 ;
        RECT 113.040 190.550 113.540 190.720 ;
        RECT 113.830 190.550 114.330 190.720 ;
        RECT 114.620 190.550 115.120 190.720 ;
        RECT 120.470 190.550 120.640 190.920 ;
        RECT 21.230 190.320 22.150 190.490 ;
        RECT 22.870 190.320 23.210 190.490 ;
        RECT 21.760 189.050 22.350 189.220 ;
        RECT 21.510 188.230 21.840 188.820 ;
        RECT 21.510 187.980 23.710 188.230 ;
        RECT 21.510 187.390 21.840 187.980 ;
        RECT 23.880 187.310 24.050 188.900 ;
        RECT 15.665 187.240 16.305 187.310 ;
        RECT 15.665 187.070 17.075 187.240 ;
        RECT 15.665 186.980 16.305 187.070 ;
        RECT 16.485 186.550 16.735 186.900 ;
        RECT 16.905 186.890 17.075 187.070 ;
        RECT 16.905 186.560 17.860 186.890 ;
        RECT 13.780 186.445 14.120 186.545 ;
        RECT 14.300 186.445 14.820 186.455 ;
        RECT 13.780 186.355 14.820 186.445 ;
        RECT 16.490 186.355 16.730 186.550 ;
        RECT 13.780 186.275 15.170 186.355 ;
        RECT 15.670 186.275 16.730 186.355 ;
        RECT 13.780 186.025 16.730 186.275 ;
        RECT 17.200 186.365 17.740 186.560 ;
        RECT 18.480 186.515 19.220 187.015 ;
        RECT 21.740 186.940 22.350 187.110 ;
        RECT 17.200 186.305 17.850 186.365 ;
        RECT 17.200 186.295 17.860 186.305 ;
        RECT 17.200 186.285 18.310 186.295 ;
        RECT 18.480 186.285 19.230 186.515 ;
        RECT 21.790 186.310 22.400 186.480 ;
        RECT 17.200 186.065 19.230 186.285 ;
        RECT 17.490 186.035 19.230 186.065 ;
        RECT 13.780 186.015 14.820 186.025 ;
        RECT 13.780 186.005 14.350 186.015 ;
        RECT 13.780 185.885 14.120 186.005 ;
        RECT 18.350 185.975 19.230 186.035 ;
        RECT 15.340 184.615 15.670 185.470 ;
        RECT 13.820 184.490 15.670 184.615 ;
        RECT 17.060 184.490 17.390 185.470 ;
        RECT 13.820 183.890 15.570 184.490 ;
        RECT 15.740 184.305 16.070 184.320 ;
        RECT 17.060 184.305 17.290 184.490 ;
        RECT 18.350 184.325 18.940 185.975 ;
        RECT 21.510 185.440 21.840 186.030 ;
        RECT 21.510 185.190 23.710 185.440 ;
        RECT 21.510 184.600 21.840 185.190 ;
        RECT 23.880 184.520 24.050 186.110 ;
        RECT 27.720 185.340 27.890 190.380 ;
        RECT 29.300 185.340 29.470 190.380 ;
        RECT 30.880 185.340 31.050 190.380 ;
        RECT 32.460 185.340 32.630 190.380 ;
        RECT 34.040 185.340 34.210 190.380 ;
        RECT 35.620 185.340 35.790 190.380 ;
        RECT 37.200 185.340 37.370 190.380 ;
        RECT 105.700 185.340 105.870 190.380 ;
        RECT 107.280 185.340 107.450 190.380 ;
        RECT 108.860 185.340 109.030 190.380 ;
        RECT 110.440 185.340 110.610 190.380 ;
        RECT 112.020 185.340 112.190 190.380 ;
        RECT 113.600 185.340 113.770 190.380 ;
        RECT 115.180 185.340 115.350 190.380 ;
        RECT 119.860 190.320 120.200 190.490 ;
        RECT 120.920 190.320 121.840 190.490 ;
        RECT 120.720 189.050 121.310 189.220 ;
        RECT 119.020 187.310 119.190 188.900 ;
        RECT 121.230 188.230 121.560 188.820 ;
        RECT 119.360 187.980 121.560 188.230 ;
        RECT 121.230 187.390 121.560 187.980 ;
        RECT 126.765 187.240 127.405 187.310 ;
        RECT 120.720 186.940 121.330 187.110 ;
        RECT 125.995 187.070 127.405 187.240 ;
        RECT 123.850 186.515 124.590 187.015 ;
        RECT 125.995 186.890 126.165 187.070 ;
        RECT 126.765 186.980 127.405 187.070 ;
        RECT 125.210 186.560 126.165 186.890 ;
        RECT 120.670 186.310 121.280 186.480 ;
        RECT 123.840 186.285 124.590 186.515 ;
        RECT 125.330 186.365 125.870 186.560 ;
        RECT 126.335 186.550 126.585 186.900 ;
        RECT 125.220 186.305 125.870 186.365 ;
        RECT 125.210 186.295 125.870 186.305 ;
        RECT 124.760 186.285 125.870 186.295 ;
        RECT 27.950 185.000 28.450 185.170 ;
        RECT 28.740 185.000 29.240 185.170 ;
        RECT 29.530 185.000 30.030 185.170 ;
        RECT 30.320 185.000 30.820 185.170 ;
        RECT 31.110 185.000 31.610 185.170 ;
        RECT 31.900 185.000 32.400 185.170 ;
        RECT 32.690 185.000 33.190 185.170 ;
        RECT 33.480 185.000 33.980 185.170 ;
        RECT 34.270 185.000 34.770 185.170 ;
        RECT 35.060 185.000 35.560 185.170 ;
        RECT 35.850 185.000 36.350 185.170 ;
        RECT 36.640 185.000 37.140 185.170 ;
        RECT 105.930 185.000 106.430 185.170 ;
        RECT 106.720 185.000 107.220 185.170 ;
        RECT 107.510 185.000 108.010 185.170 ;
        RECT 108.300 185.000 108.800 185.170 ;
        RECT 109.090 185.000 109.590 185.170 ;
        RECT 109.880 185.000 110.380 185.170 ;
        RECT 110.670 185.000 111.170 185.170 ;
        RECT 111.460 185.000 111.960 185.170 ;
        RECT 112.250 185.000 112.750 185.170 ;
        RECT 113.040 185.000 113.540 185.170 ;
        RECT 113.830 185.000 114.330 185.170 ;
        RECT 114.620 185.000 115.120 185.170 ;
        RECT 119.020 184.520 119.190 186.110 ;
        RECT 123.840 186.065 125.870 186.285 ;
        RECT 126.340 186.355 126.580 186.550 ;
        RECT 128.250 186.445 128.770 186.455 ;
        RECT 128.950 186.445 129.290 186.545 ;
        RECT 128.250 186.355 129.290 186.445 ;
        RECT 126.340 186.275 127.400 186.355 ;
        RECT 127.900 186.275 129.290 186.355 ;
        RECT 123.840 186.035 125.580 186.065 ;
        RECT 121.230 185.440 121.560 186.030 ;
        RECT 123.840 185.975 124.720 186.035 ;
        RECT 126.340 186.025 129.290 186.275 ;
        RECT 128.250 186.015 129.290 186.025 ;
        RECT 128.720 186.005 129.290 186.015 ;
        RECT 119.360 185.190 121.560 185.440 ;
        RECT 121.230 184.600 121.560 185.190 ;
        RECT 17.580 184.320 18.940 184.325 ;
        RECT 15.740 184.085 17.290 184.305 ;
        RECT 15.740 184.080 16.070 184.085 ;
        RECT 17.060 183.890 17.290 184.085 ;
        RECT 17.460 184.085 18.940 184.320 ;
        RECT 21.760 184.200 22.350 184.370 ;
        RECT 120.720 184.200 121.310 184.370 ;
        RECT 124.130 184.325 124.720 185.975 ;
        RECT 128.950 185.885 129.290 186.005 ;
        RECT 125.680 184.490 126.010 185.470 ;
        RECT 127.400 184.615 127.730 185.470 ;
        RECT 127.400 184.490 129.250 184.615 ;
        RECT 124.130 184.320 125.490 184.325 ;
        RECT 124.130 184.085 125.610 184.320 ;
        RECT 17.460 184.080 17.790 184.085 ;
        RECT 125.280 184.080 125.610 184.085 ;
        RECT 125.780 184.305 126.010 184.490 ;
        RECT 127.000 184.305 127.330 184.320 ;
        RECT 125.780 184.085 127.330 184.305 ;
        RECT 125.780 183.890 126.010 184.085 ;
        RECT 127.000 184.080 127.330 184.085 ;
        RECT 127.500 183.890 129.250 184.490 ;
        RECT 13.820 183.825 15.670 183.890 ;
        RECT 15.340 183.260 15.670 183.825 ;
        RECT 17.060 183.260 17.390 183.890 ;
        RECT 125.680 183.260 126.010 183.890 ;
        RECT 127.400 183.825 129.250 183.890 ;
        RECT 127.400 183.260 127.730 183.825 ;
        RECT 23.060 182.070 23.560 182.240 ;
        RECT 23.850 182.070 24.350 182.240 ;
        RECT 24.640 182.070 25.140 182.240 ;
        RECT 25.430 182.070 25.930 182.240 ;
        RECT 26.220 182.070 26.720 182.240 ;
        RECT 27.010 182.070 27.510 182.240 ;
        RECT 27.800 182.070 28.300 182.240 ;
        RECT 28.590 182.070 29.090 182.240 ;
        RECT 29.380 182.070 29.880 182.240 ;
        RECT 30.170 182.070 30.670 182.240 ;
        RECT 30.960 182.070 31.460 182.240 ;
        RECT 31.750 182.070 32.250 182.240 ;
        RECT 32.540 182.070 33.040 182.240 ;
        RECT 33.330 182.070 33.830 182.240 ;
        RECT 34.120 182.070 34.620 182.240 ;
        RECT 34.910 182.070 35.410 182.240 ;
        RECT 35.700 182.070 36.200 182.240 ;
        RECT 36.490 182.070 36.990 182.240 ;
        RECT 106.080 182.070 106.580 182.240 ;
        RECT 106.870 182.070 107.370 182.240 ;
        RECT 107.660 182.070 108.160 182.240 ;
        RECT 108.450 182.070 108.950 182.240 ;
        RECT 109.240 182.070 109.740 182.240 ;
        RECT 110.030 182.070 110.530 182.240 ;
        RECT 110.820 182.070 111.320 182.240 ;
        RECT 111.610 182.070 112.110 182.240 ;
        RECT 112.400 182.070 112.900 182.240 ;
        RECT 113.190 182.070 113.690 182.240 ;
        RECT 113.980 182.070 114.480 182.240 ;
        RECT 114.770 182.070 115.270 182.240 ;
        RECT 115.560 182.070 116.060 182.240 ;
        RECT 116.350 182.070 116.850 182.240 ;
        RECT 117.140 182.070 117.640 182.240 ;
        RECT 117.930 182.070 118.430 182.240 ;
        RECT 118.720 182.070 119.220 182.240 ;
        RECT 119.510 182.070 120.010 182.240 ;
        RECT 15.500 181.135 15.830 181.360 ;
        RECT 15.120 180.575 15.830 181.135 ;
        RECT 15.500 180.380 15.830 180.575 ;
        RECT 17.160 180.390 17.490 181.370 ;
        RECT 15.500 179.780 15.730 180.380 ;
        RECT 15.900 180.175 16.230 180.210 ;
        RECT 17.160 180.175 17.390 180.390 ;
        RECT 15.900 179.985 17.390 180.175 ;
        RECT 15.900 179.970 16.230 179.985 ;
        RECT 17.160 179.790 17.390 179.985 ;
        RECT 17.560 180.215 17.890 180.220 ;
        RECT 18.200 180.215 19.030 180.305 ;
        RECT 17.560 179.985 19.030 180.215 ;
        RECT 17.560 179.980 17.890 179.985 ;
        RECT 15.500 179.150 15.830 179.780 ;
        RECT 17.160 179.160 17.490 179.790 ;
        RECT 18.200 179.785 19.030 179.985 ;
        RECT 14.580 178.245 16.660 178.565 ;
        RECT 14.580 178.165 15.100 178.245 ;
        RECT 15.590 178.165 16.660 178.245 ;
        RECT 16.420 177.990 16.660 178.165 ;
        RECT 16.415 177.640 16.665 177.990 ;
        RECT 15.595 177.470 16.235 177.540 ;
        RECT 15.595 177.300 17.005 177.470 ;
        RECT 15.595 177.210 16.235 177.300 ;
        RECT 16.415 176.780 16.665 177.130 ;
        RECT 16.835 177.120 17.005 177.300 ;
        RECT 16.835 176.790 17.790 177.120 ;
        RECT 16.420 176.605 16.660 176.780 ;
        RECT 16.420 176.145 16.670 176.605 ;
        RECT 15.565 175.915 17.775 176.145 ;
        RECT 15.565 175.815 16.195 175.915 ;
        RECT 16.795 175.815 17.775 175.915 ;
        RECT 22.830 171.815 23.000 181.855 ;
        RECT 24.410 171.815 24.580 181.855 ;
        RECT 25.990 171.815 26.160 181.855 ;
        RECT 27.570 171.815 27.740 181.855 ;
        RECT 29.150 171.815 29.320 181.855 ;
        RECT 30.730 171.815 30.900 181.855 ;
        RECT 32.310 171.815 32.480 181.855 ;
        RECT 33.890 171.815 34.060 181.855 ;
        RECT 35.470 171.815 35.640 181.855 ;
        RECT 37.050 171.815 37.220 181.855 ;
        RECT 105.850 171.815 106.020 181.855 ;
        RECT 107.430 171.815 107.600 181.855 ;
        RECT 109.010 171.815 109.180 181.855 ;
        RECT 110.590 171.815 110.760 181.855 ;
        RECT 112.170 171.815 112.340 181.855 ;
        RECT 113.750 171.815 113.920 181.855 ;
        RECT 115.330 171.815 115.500 181.855 ;
        RECT 116.910 171.815 117.080 181.855 ;
        RECT 118.490 171.815 118.660 181.855 ;
        RECT 120.070 171.815 120.240 181.855 ;
        RECT 125.580 180.390 125.910 181.370 ;
        RECT 124.040 180.215 124.870 180.305 ;
        RECT 125.180 180.215 125.510 180.220 ;
        RECT 124.040 179.985 125.510 180.215 ;
        RECT 124.040 179.785 124.870 179.985 ;
        RECT 125.180 179.980 125.510 179.985 ;
        RECT 125.680 180.175 125.910 180.390 ;
        RECT 127.240 181.135 127.570 181.360 ;
        RECT 127.240 180.575 127.950 181.135 ;
        RECT 127.240 180.380 127.570 180.575 ;
        RECT 126.840 180.175 127.170 180.210 ;
        RECT 125.680 179.985 127.170 180.175 ;
        RECT 125.680 179.790 125.910 179.985 ;
        RECT 126.840 179.970 127.170 179.985 ;
        RECT 125.580 179.160 125.910 179.790 ;
        RECT 127.340 179.780 127.570 180.380 ;
        RECT 127.240 179.150 127.570 179.780 ;
        RECT 126.410 178.245 128.490 178.565 ;
        RECT 126.410 178.165 127.480 178.245 ;
        RECT 127.970 178.165 128.490 178.245 ;
        RECT 126.410 177.990 126.650 178.165 ;
        RECT 126.405 177.640 126.655 177.990 ;
        RECT 126.835 177.470 127.475 177.540 ;
        RECT 126.065 177.300 127.475 177.470 ;
        RECT 126.065 177.120 126.235 177.300 ;
        RECT 126.835 177.210 127.475 177.300 ;
        RECT 125.280 176.790 126.235 177.120 ;
        RECT 126.405 176.780 126.655 177.130 ;
        RECT 126.410 176.605 126.650 176.780 ;
        RECT 126.400 176.145 126.650 176.605 ;
        RECT 125.295 175.915 127.505 176.145 ;
        RECT 125.295 175.815 126.275 175.915 ;
        RECT 126.875 175.815 127.505 175.915 ;
        RECT 23.060 171.430 23.560 171.600 ;
        RECT 23.850 171.430 24.350 171.600 ;
        RECT 24.640 171.430 25.140 171.600 ;
        RECT 25.430 171.430 25.930 171.600 ;
        RECT 26.220 171.430 26.720 171.600 ;
        RECT 27.010 171.430 27.510 171.600 ;
        RECT 27.800 171.430 28.300 171.600 ;
        RECT 28.590 171.430 29.090 171.600 ;
        RECT 29.380 171.430 29.880 171.600 ;
        RECT 30.170 171.430 30.670 171.600 ;
        RECT 30.960 171.430 31.460 171.600 ;
        RECT 31.750 171.430 32.250 171.600 ;
        RECT 32.540 171.430 33.040 171.600 ;
        RECT 33.330 171.430 33.830 171.600 ;
        RECT 34.120 171.430 34.620 171.600 ;
        RECT 34.910 171.430 35.410 171.600 ;
        RECT 35.700 171.430 36.200 171.600 ;
        RECT 36.490 171.430 36.990 171.600 ;
        RECT 106.080 171.430 106.580 171.600 ;
        RECT 106.870 171.430 107.370 171.600 ;
        RECT 107.660 171.430 108.160 171.600 ;
        RECT 108.450 171.430 108.950 171.600 ;
        RECT 109.240 171.430 109.740 171.600 ;
        RECT 110.030 171.430 110.530 171.600 ;
        RECT 110.820 171.430 111.320 171.600 ;
        RECT 111.610 171.430 112.110 171.600 ;
        RECT 112.400 171.430 112.900 171.600 ;
        RECT 113.190 171.430 113.690 171.600 ;
        RECT 113.980 171.430 114.480 171.600 ;
        RECT 114.770 171.430 115.270 171.600 ;
        RECT 115.560 171.430 116.060 171.600 ;
        RECT 116.350 171.430 116.850 171.600 ;
        RECT 117.140 171.430 117.640 171.600 ;
        RECT 117.930 171.430 118.430 171.600 ;
        RECT 118.720 171.430 119.220 171.600 ;
        RECT 119.510 171.430 120.010 171.600 ;
        RECT 22.905 165.295 23.405 165.465 ;
        RECT 23.695 165.295 24.195 165.465 ;
        RECT 24.485 165.295 24.985 165.465 ;
        RECT 25.275 165.295 25.775 165.465 ;
        RECT 26.065 165.295 26.565 165.465 ;
        RECT 26.855 165.295 27.355 165.465 ;
        RECT 27.645 165.295 28.145 165.465 ;
        RECT 28.435 165.295 28.935 165.465 ;
        RECT 29.225 165.295 29.725 165.465 ;
        RECT 30.015 165.295 30.515 165.465 ;
        RECT 30.805 165.295 31.305 165.465 ;
        RECT 31.595 165.295 32.095 165.465 ;
        RECT 32.385 165.295 32.885 165.465 ;
        RECT 33.175 165.295 33.675 165.465 ;
        RECT 33.965 165.295 34.465 165.465 ;
        RECT 34.755 165.295 35.255 165.465 ;
        RECT 35.545 165.295 36.045 165.465 ;
        RECT 36.335 165.295 36.835 165.465 ;
        RECT 106.235 165.295 106.735 165.465 ;
        RECT 107.025 165.295 107.525 165.465 ;
        RECT 107.815 165.295 108.315 165.465 ;
        RECT 108.605 165.295 109.105 165.465 ;
        RECT 109.395 165.295 109.895 165.465 ;
        RECT 110.185 165.295 110.685 165.465 ;
        RECT 110.975 165.295 111.475 165.465 ;
        RECT 111.765 165.295 112.265 165.465 ;
        RECT 112.555 165.295 113.055 165.465 ;
        RECT 113.345 165.295 113.845 165.465 ;
        RECT 114.135 165.295 114.635 165.465 ;
        RECT 114.925 165.295 115.425 165.465 ;
        RECT 115.715 165.295 116.215 165.465 ;
        RECT 116.505 165.295 117.005 165.465 ;
        RECT 117.295 165.295 117.795 165.465 ;
        RECT 118.085 165.295 118.585 165.465 ;
        RECT 118.875 165.295 119.375 165.465 ;
        RECT 119.665 165.295 120.165 165.465 ;
        RECT 22.675 155.040 22.845 165.080 ;
        RECT 24.255 155.040 24.425 165.080 ;
        RECT 25.835 155.040 26.005 165.080 ;
        RECT 27.415 155.040 27.585 165.080 ;
        RECT 28.995 155.040 29.165 165.080 ;
        RECT 30.575 155.040 30.745 165.080 ;
        RECT 32.155 155.040 32.325 165.080 ;
        RECT 33.735 155.040 33.905 165.080 ;
        RECT 35.315 155.040 35.485 165.080 ;
        RECT 36.895 155.040 37.065 165.080 ;
        RECT 106.005 155.040 106.175 165.080 ;
        RECT 107.585 155.040 107.755 165.080 ;
        RECT 109.165 155.040 109.335 165.080 ;
        RECT 110.745 155.040 110.915 165.080 ;
        RECT 112.325 155.040 112.495 165.080 ;
        RECT 113.905 155.040 114.075 165.080 ;
        RECT 115.485 155.040 115.655 165.080 ;
        RECT 117.065 155.040 117.235 165.080 ;
        RECT 118.645 155.040 118.815 165.080 ;
        RECT 120.225 155.040 120.395 165.080 ;
        RECT 22.905 154.655 23.405 154.825 ;
        RECT 23.695 154.655 24.195 154.825 ;
        RECT 24.485 154.655 24.985 154.825 ;
        RECT 25.275 154.655 25.775 154.825 ;
        RECT 26.065 154.655 26.565 154.825 ;
        RECT 26.855 154.655 27.355 154.825 ;
        RECT 27.645 154.655 28.145 154.825 ;
        RECT 28.435 154.655 28.935 154.825 ;
        RECT 29.225 154.655 29.725 154.825 ;
        RECT 30.015 154.655 30.515 154.825 ;
        RECT 30.805 154.655 31.305 154.825 ;
        RECT 31.595 154.655 32.095 154.825 ;
        RECT 32.385 154.655 32.885 154.825 ;
        RECT 33.175 154.655 33.675 154.825 ;
        RECT 33.965 154.655 34.465 154.825 ;
        RECT 34.755 154.655 35.255 154.825 ;
        RECT 35.545 154.655 36.045 154.825 ;
        RECT 36.335 154.655 36.835 154.825 ;
        RECT 106.235 154.655 106.735 154.825 ;
        RECT 107.025 154.655 107.525 154.825 ;
        RECT 107.815 154.655 108.315 154.825 ;
        RECT 108.605 154.655 109.105 154.825 ;
        RECT 109.395 154.655 109.895 154.825 ;
        RECT 110.185 154.655 110.685 154.825 ;
        RECT 110.975 154.655 111.475 154.825 ;
        RECT 111.765 154.655 112.265 154.825 ;
        RECT 112.555 154.655 113.055 154.825 ;
        RECT 113.345 154.655 113.845 154.825 ;
        RECT 114.135 154.655 114.635 154.825 ;
        RECT 114.925 154.655 115.425 154.825 ;
        RECT 115.715 154.655 116.215 154.825 ;
        RECT 116.505 154.655 117.005 154.825 ;
        RECT 117.295 154.655 117.795 154.825 ;
        RECT 118.085 154.655 118.585 154.825 ;
        RECT 118.875 154.655 119.375 154.825 ;
        RECT 119.665 154.655 120.165 154.825 ;
        RECT 37.545 152.525 38.135 152.695 ;
        RECT 104.935 152.525 105.525 152.695 ;
        RECT 22.755 151.725 23.255 151.895 ;
        RECT 23.545 151.725 24.045 151.895 ;
        RECT 24.335 151.725 24.835 151.895 ;
        RECT 25.125 151.725 25.625 151.895 ;
        RECT 25.915 151.725 26.415 151.895 ;
        RECT 26.705 151.725 27.205 151.895 ;
        RECT 27.495 151.725 27.995 151.895 ;
        RECT 28.285 151.725 28.785 151.895 ;
        RECT 29.075 151.725 29.575 151.895 ;
        RECT 29.865 151.725 30.365 151.895 ;
        RECT 30.655 151.725 31.155 151.895 ;
        RECT 31.445 151.725 31.945 151.895 ;
        RECT 22.525 146.515 22.695 151.555 ;
        RECT 24.105 146.515 24.275 151.555 ;
        RECT 25.685 146.515 25.855 151.555 ;
        RECT 27.265 146.515 27.435 151.555 ;
        RECT 28.845 146.515 29.015 151.555 ;
        RECT 30.425 146.515 30.595 151.555 ;
        RECT 32.005 146.515 32.175 151.555 ;
        RECT 35.845 150.785 36.015 152.375 ;
        RECT 38.055 151.705 38.385 152.295 ;
        RECT 36.185 151.455 38.385 151.705 ;
        RECT 38.055 150.865 38.385 151.455 ;
        RECT 104.685 151.705 105.015 152.295 ;
        RECT 104.685 151.455 106.885 151.705 ;
        RECT 104.685 150.865 105.015 151.455 ;
        RECT 107.055 150.785 107.225 152.375 ;
        RECT 111.125 151.725 111.625 151.895 ;
        RECT 111.915 151.725 112.415 151.895 ;
        RECT 112.705 151.725 113.205 151.895 ;
        RECT 113.495 151.725 113.995 151.895 ;
        RECT 114.285 151.725 114.785 151.895 ;
        RECT 115.075 151.725 115.575 151.895 ;
        RECT 115.865 151.725 116.365 151.895 ;
        RECT 116.655 151.725 117.155 151.895 ;
        RECT 117.445 151.725 117.945 151.895 ;
        RECT 118.235 151.725 118.735 151.895 ;
        RECT 119.025 151.725 119.525 151.895 ;
        RECT 119.815 151.725 120.315 151.895 ;
        RECT 37.495 150.415 38.105 150.585 ;
        RECT 104.965 150.415 105.575 150.585 ;
        RECT 37.545 149.785 38.155 149.955 ;
        RECT 104.915 149.785 105.525 149.955 ;
        RECT 35.845 147.995 36.015 149.585 ;
        RECT 38.055 148.915 38.385 149.505 ;
        RECT 36.185 148.665 38.385 148.915 ;
        RECT 38.055 148.075 38.385 148.665 ;
        RECT 104.685 148.915 105.015 149.505 ;
        RECT 104.685 148.665 106.885 148.915 ;
        RECT 104.685 148.075 105.015 148.665 ;
        RECT 107.055 147.995 107.225 149.585 ;
        RECT 37.545 147.675 38.135 147.845 ;
        RECT 104.935 147.675 105.525 147.845 ;
        RECT 36.685 146.405 37.025 146.575 ;
        RECT 37.745 146.405 38.665 146.575 ;
        RECT 104.405 146.405 105.325 146.575 ;
        RECT 106.045 146.405 106.385 146.575 ;
        RECT 110.895 146.515 111.065 151.555 ;
        RECT 112.475 146.515 112.645 151.555 ;
        RECT 114.055 146.515 114.225 151.555 ;
        RECT 115.635 146.515 115.805 151.555 ;
        RECT 117.215 146.515 117.385 151.555 ;
        RECT 118.795 146.515 118.965 151.555 ;
        RECT 120.375 146.515 120.545 151.555 ;
        RECT 22.755 146.175 23.255 146.345 ;
        RECT 23.545 146.175 24.045 146.345 ;
        RECT 24.335 146.175 24.835 146.345 ;
        RECT 25.125 146.175 25.625 146.345 ;
        RECT 25.915 146.175 26.415 146.345 ;
        RECT 26.705 146.175 27.205 146.345 ;
        RECT 27.495 146.175 27.995 146.345 ;
        RECT 28.285 146.175 28.785 146.345 ;
        RECT 29.075 146.175 29.575 146.345 ;
        RECT 29.865 146.175 30.365 146.345 ;
        RECT 30.655 146.175 31.155 146.345 ;
        RECT 31.445 146.175 31.945 146.345 ;
        RECT 37.295 145.975 37.465 146.345 ;
        RECT 105.605 145.975 105.775 146.345 ;
        RECT 111.125 146.175 111.625 146.345 ;
        RECT 111.915 146.175 112.415 146.345 ;
        RECT 112.705 146.175 113.205 146.345 ;
        RECT 113.495 146.175 113.995 146.345 ;
        RECT 114.285 146.175 114.785 146.345 ;
        RECT 115.075 146.175 115.575 146.345 ;
        RECT 115.865 146.175 116.365 146.345 ;
        RECT 116.655 146.175 117.155 146.345 ;
        RECT 117.445 146.175 117.945 146.345 ;
        RECT 118.235 146.175 118.735 146.345 ;
        RECT 119.025 146.175 119.525 146.345 ;
        RECT 119.815 146.175 120.315 146.345 ;
        RECT 22.430 140.980 22.600 141.350 ;
        RECT 27.950 140.980 28.450 141.150 ;
        RECT 28.740 140.980 29.240 141.150 ;
        RECT 29.530 140.980 30.030 141.150 ;
        RECT 30.320 140.980 30.820 141.150 ;
        RECT 31.110 140.980 31.610 141.150 ;
        RECT 31.900 140.980 32.400 141.150 ;
        RECT 32.690 140.980 33.190 141.150 ;
        RECT 33.480 140.980 33.980 141.150 ;
        RECT 34.270 140.980 34.770 141.150 ;
        RECT 35.060 140.980 35.560 141.150 ;
        RECT 35.850 140.980 36.350 141.150 ;
        RECT 36.640 140.980 37.140 141.150 ;
        RECT 105.930 140.980 106.430 141.150 ;
        RECT 106.720 140.980 107.220 141.150 ;
        RECT 107.510 140.980 108.010 141.150 ;
        RECT 108.300 140.980 108.800 141.150 ;
        RECT 109.090 140.980 109.590 141.150 ;
        RECT 109.880 140.980 110.380 141.150 ;
        RECT 110.670 140.980 111.170 141.150 ;
        RECT 111.460 140.980 111.960 141.150 ;
        RECT 112.250 140.980 112.750 141.150 ;
        RECT 113.040 140.980 113.540 141.150 ;
        RECT 113.830 140.980 114.330 141.150 ;
        RECT 114.620 140.980 115.120 141.150 ;
        RECT 120.470 140.980 120.640 141.350 ;
        RECT 21.230 140.750 22.150 140.920 ;
        RECT 22.870 140.750 23.210 140.920 ;
        RECT 21.760 139.480 22.350 139.650 ;
        RECT 21.510 138.660 21.840 139.250 ;
        RECT 21.510 138.410 23.710 138.660 ;
        RECT 21.510 137.820 21.840 138.410 ;
        RECT 23.880 137.740 24.050 139.330 ;
        RECT 15.665 137.670 16.305 137.740 ;
        RECT 15.665 137.500 17.075 137.670 ;
        RECT 15.665 137.410 16.305 137.500 ;
        RECT 16.485 136.980 16.735 137.330 ;
        RECT 16.905 137.320 17.075 137.500 ;
        RECT 16.905 136.990 17.860 137.320 ;
        RECT 13.780 136.875 14.120 136.975 ;
        RECT 14.300 136.875 14.820 136.885 ;
        RECT 13.780 136.785 14.820 136.875 ;
        RECT 16.490 136.785 16.730 136.980 ;
        RECT 13.780 136.705 15.170 136.785 ;
        RECT 15.670 136.705 16.730 136.785 ;
        RECT 13.780 136.455 16.730 136.705 ;
        RECT 17.200 136.795 17.740 136.990 ;
        RECT 18.480 136.945 19.220 137.445 ;
        RECT 21.740 137.370 22.350 137.540 ;
        RECT 17.200 136.735 17.850 136.795 ;
        RECT 17.200 136.725 17.860 136.735 ;
        RECT 17.200 136.715 18.310 136.725 ;
        RECT 18.480 136.715 19.230 136.945 ;
        RECT 21.790 136.740 22.400 136.910 ;
        RECT 17.200 136.495 19.230 136.715 ;
        RECT 17.490 136.465 19.230 136.495 ;
        RECT 13.780 136.445 14.820 136.455 ;
        RECT 13.780 136.435 14.350 136.445 ;
        RECT 13.780 136.315 14.120 136.435 ;
        RECT 18.350 136.405 19.230 136.465 ;
        RECT 15.340 135.045 15.670 135.900 ;
        RECT 13.820 134.920 15.670 135.045 ;
        RECT 17.060 134.920 17.390 135.900 ;
        RECT 13.820 134.320 15.570 134.920 ;
        RECT 15.740 134.735 16.070 134.750 ;
        RECT 17.060 134.735 17.290 134.920 ;
        RECT 18.350 134.755 18.940 136.405 ;
        RECT 21.510 135.870 21.840 136.460 ;
        RECT 21.510 135.620 23.710 135.870 ;
        RECT 21.510 135.030 21.840 135.620 ;
        RECT 23.880 134.950 24.050 136.540 ;
        RECT 27.720 135.770 27.890 140.810 ;
        RECT 29.300 135.770 29.470 140.810 ;
        RECT 30.880 135.770 31.050 140.810 ;
        RECT 32.460 135.770 32.630 140.810 ;
        RECT 34.040 135.770 34.210 140.810 ;
        RECT 35.620 135.770 35.790 140.810 ;
        RECT 37.200 135.770 37.370 140.810 ;
        RECT 105.700 135.770 105.870 140.810 ;
        RECT 107.280 135.770 107.450 140.810 ;
        RECT 108.860 135.770 109.030 140.810 ;
        RECT 110.440 135.770 110.610 140.810 ;
        RECT 112.020 135.770 112.190 140.810 ;
        RECT 113.600 135.770 113.770 140.810 ;
        RECT 115.180 135.770 115.350 140.810 ;
        RECT 119.860 140.750 120.200 140.920 ;
        RECT 120.920 140.750 121.840 140.920 ;
        RECT 120.720 139.480 121.310 139.650 ;
        RECT 119.020 137.740 119.190 139.330 ;
        RECT 121.230 138.660 121.560 139.250 ;
        RECT 119.360 138.410 121.560 138.660 ;
        RECT 121.230 137.820 121.560 138.410 ;
        RECT 126.765 137.670 127.405 137.740 ;
        RECT 120.720 137.370 121.330 137.540 ;
        RECT 125.995 137.500 127.405 137.670 ;
        RECT 123.850 136.945 124.590 137.445 ;
        RECT 125.995 137.320 126.165 137.500 ;
        RECT 126.765 137.410 127.405 137.500 ;
        RECT 125.210 136.990 126.165 137.320 ;
        RECT 120.670 136.740 121.280 136.910 ;
        RECT 123.840 136.715 124.590 136.945 ;
        RECT 125.330 136.795 125.870 136.990 ;
        RECT 126.335 136.980 126.585 137.330 ;
        RECT 125.220 136.735 125.870 136.795 ;
        RECT 125.210 136.725 125.870 136.735 ;
        RECT 124.760 136.715 125.870 136.725 ;
        RECT 27.950 135.430 28.450 135.600 ;
        RECT 28.740 135.430 29.240 135.600 ;
        RECT 29.530 135.430 30.030 135.600 ;
        RECT 30.320 135.430 30.820 135.600 ;
        RECT 31.110 135.430 31.610 135.600 ;
        RECT 31.900 135.430 32.400 135.600 ;
        RECT 32.690 135.430 33.190 135.600 ;
        RECT 33.480 135.430 33.980 135.600 ;
        RECT 34.270 135.430 34.770 135.600 ;
        RECT 35.060 135.430 35.560 135.600 ;
        RECT 35.850 135.430 36.350 135.600 ;
        RECT 36.640 135.430 37.140 135.600 ;
        RECT 105.930 135.430 106.430 135.600 ;
        RECT 106.720 135.430 107.220 135.600 ;
        RECT 107.510 135.430 108.010 135.600 ;
        RECT 108.300 135.430 108.800 135.600 ;
        RECT 109.090 135.430 109.590 135.600 ;
        RECT 109.880 135.430 110.380 135.600 ;
        RECT 110.670 135.430 111.170 135.600 ;
        RECT 111.460 135.430 111.960 135.600 ;
        RECT 112.250 135.430 112.750 135.600 ;
        RECT 113.040 135.430 113.540 135.600 ;
        RECT 113.830 135.430 114.330 135.600 ;
        RECT 114.620 135.430 115.120 135.600 ;
        RECT 119.020 134.950 119.190 136.540 ;
        RECT 123.840 136.495 125.870 136.715 ;
        RECT 126.340 136.785 126.580 136.980 ;
        RECT 128.250 136.875 128.770 136.885 ;
        RECT 128.950 136.875 129.290 136.975 ;
        RECT 128.250 136.785 129.290 136.875 ;
        RECT 126.340 136.705 127.400 136.785 ;
        RECT 127.900 136.705 129.290 136.785 ;
        RECT 123.840 136.465 125.580 136.495 ;
        RECT 121.230 135.870 121.560 136.460 ;
        RECT 123.840 136.405 124.720 136.465 ;
        RECT 126.340 136.455 129.290 136.705 ;
        RECT 128.250 136.445 129.290 136.455 ;
        RECT 128.720 136.435 129.290 136.445 ;
        RECT 119.360 135.620 121.560 135.870 ;
        RECT 121.230 135.030 121.560 135.620 ;
        RECT 17.580 134.750 18.940 134.755 ;
        RECT 15.740 134.515 17.290 134.735 ;
        RECT 15.740 134.510 16.070 134.515 ;
        RECT 17.060 134.320 17.290 134.515 ;
        RECT 17.460 134.515 18.940 134.750 ;
        RECT 21.760 134.630 22.350 134.800 ;
        RECT 120.720 134.630 121.310 134.800 ;
        RECT 124.130 134.755 124.720 136.405 ;
        RECT 128.950 136.315 129.290 136.435 ;
        RECT 125.680 134.920 126.010 135.900 ;
        RECT 127.400 135.045 127.730 135.900 ;
        RECT 127.400 134.920 129.250 135.045 ;
        RECT 124.130 134.750 125.490 134.755 ;
        RECT 124.130 134.515 125.610 134.750 ;
        RECT 17.460 134.510 17.790 134.515 ;
        RECT 125.280 134.510 125.610 134.515 ;
        RECT 125.780 134.735 126.010 134.920 ;
        RECT 127.000 134.735 127.330 134.750 ;
        RECT 125.780 134.515 127.330 134.735 ;
        RECT 125.780 134.320 126.010 134.515 ;
        RECT 127.000 134.510 127.330 134.515 ;
        RECT 127.500 134.320 129.250 134.920 ;
        RECT 13.820 134.255 15.670 134.320 ;
        RECT 15.340 133.690 15.670 134.255 ;
        RECT 17.060 133.690 17.390 134.320 ;
        RECT 125.680 133.690 126.010 134.320 ;
        RECT 127.400 134.255 129.250 134.320 ;
        RECT 127.400 133.690 127.730 134.255 ;
        RECT 23.060 132.500 23.560 132.670 ;
        RECT 23.850 132.500 24.350 132.670 ;
        RECT 24.640 132.500 25.140 132.670 ;
        RECT 25.430 132.500 25.930 132.670 ;
        RECT 26.220 132.500 26.720 132.670 ;
        RECT 27.010 132.500 27.510 132.670 ;
        RECT 27.800 132.500 28.300 132.670 ;
        RECT 28.590 132.500 29.090 132.670 ;
        RECT 29.380 132.500 29.880 132.670 ;
        RECT 30.170 132.500 30.670 132.670 ;
        RECT 30.960 132.500 31.460 132.670 ;
        RECT 31.750 132.500 32.250 132.670 ;
        RECT 32.540 132.500 33.040 132.670 ;
        RECT 33.330 132.500 33.830 132.670 ;
        RECT 34.120 132.500 34.620 132.670 ;
        RECT 34.910 132.500 35.410 132.670 ;
        RECT 35.700 132.500 36.200 132.670 ;
        RECT 36.490 132.500 36.990 132.670 ;
        RECT 106.080 132.500 106.580 132.670 ;
        RECT 106.870 132.500 107.370 132.670 ;
        RECT 107.660 132.500 108.160 132.670 ;
        RECT 108.450 132.500 108.950 132.670 ;
        RECT 109.240 132.500 109.740 132.670 ;
        RECT 110.030 132.500 110.530 132.670 ;
        RECT 110.820 132.500 111.320 132.670 ;
        RECT 111.610 132.500 112.110 132.670 ;
        RECT 112.400 132.500 112.900 132.670 ;
        RECT 113.190 132.500 113.690 132.670 ;
        RECT 113.980 132.500 114.480 132.670 ;
        RECT 114.770 132.500 115.270 132.670 ;
        RECT 115.560 132.500 116.060 132.670 ;
        RECT 116.350 132.500 116.850 132.670 ;
        RECT 117.140 132.500 117.640 132.670 ;
        RECT 117.930 132.500 118.430 132.670 ;
        RECT 118.720 132.500 119.220 132.670 ;
        RECT 119.510 132.500 120.010 132.670 ;
        RECT 15.500 131.565 15.830 131.790 ;
        RECT 15.120 131.005 15.830 131.565 ;
        RECT 15.500 130.810 15.830 131.005 ;
        RECT 17.160 130.820 17.490 131.800 ;
        RECT 15.500 130.210 15.730 130.810 ;
        RECT 15.900 130.605 16.230 130.640 ;
        RECT 17.160 130.605 17.390 130.820 ;
        RECT 15.900 130.415 17.390 130.605 ;
        RECT 15.900 130.400 16.230 130.415 ;
        RECT 17.160 130.220 17.390 130.415 ;
        RECT 17.560 130.645 17.890 130.650 ;
        RECT 18.200 130.645 19.030 130.735 ;
        RECT 17.560 130.415 19.030 130.645 ;
        RECT 17.560 130.410 17.890 130.415 ;
        RECT 15.500 129.580 15.830 130.210 ;
        RECT 17.160 129.590 17.490 130.220 ;
        RECT 18.200 130.215 19.030 130.415 ;
        RECT 14.580 128.675 16.660 128.995 ;
        RECT 14.580 128.595 15.100 128.675 ;
        RECT 15.590 128.595 16.660 128.675 ;
        RECT 16.420 128.420 16.660 128.595 ;
        RECT 16.415 128.070 16.665 128.420 ;
        RECT 15.595 127.900 16.235 127.970 ;
        RECT 15.595 127.730 17.005 127.900 ;
        RECT 15.595 127.640 16.235 127.730 ;
        RECT 16.415 127.210 16.665 127.560 ;
        RECT 16.835 127.550 17.005 127.730 ;
        RECT 16.835 127.220 17.790 127.550 ;
        RECT 16.420 127.035 16.660 127.210 ;
        RECT 16.420 126.575 16.670 127.035 ;
        RECT 15.565 126.345 17.775 126.575 ;
        RECT 15.565 126.245 16.195 126.345 ;
        RECT 16.795 126.245 17.775 126.345 ;
        RECT 22.830 122.245 23.000 132.285 ;
        RECT 24.410 122.245 24.580 132.285 ;
        RECT 25.990 122.245 26.160 132.285 ;
        RECT 27.570 122.245 27.740 132.285 ;
        RECT 29.150 122.245 29.320 132.285 ;
        RECT 30.730 122.245 30.900 132.285 ;
        RECT 32.310 122.245 32.480 132.285 ;
        RECT 33.890 122.245 34.060 132.285 ;
        RECT 35.470 122.245 35.640 132.285 ;
        RECT 37.050 122.245 37.220 132.285 ;
        RECT 105.850 122.245 106.020 132.285 ;
        RECT 107.430 122.245 107.600 132.285 ;
        RECT 109.010 122.245 109.180 132.285 ;
        RECT 110.590 122.245 110.760 132.285 ;
        RECT 112.170 122.245 112.340 132.285 ;
        RECT 113.750 122.245 113.920 132.285 ;
        RECT 115.330 122.245 115.500 132.285 ;
        RECT 116.910 122.245 117.080 132.285 ;
        RECT 118.490 122.245 118.660 132.285 ;
        RECT 120.070 122.245 120.240 132.285 ;
        RECT 125.580 130.820 125.910 131.800 ;
        RECT 124.040 130.645 124.870 130.735 ;
        RECT 125.180 130.645 125.510 130.650 ;
        RECT 124.040 130.415 125.510 130.645 ;
        RECT 124.040 130.215 124.870 130.415 ;
        RECT 125.180 130.410 125.510 130.415 ;
        RECT 125.680 130.605 125.910 130.820 ;
        RECT 127.240 131.565 127.570 131.790 ;
        RECT 127.240 131.005 127.950 131.565 ;
        RECT 127.240 130.810 127.570 131.005 ;
        RECT 126.840 130.605 127.170 130.640 ;
        RECT 125.680 130.415 127.170 130.605 ;
        RECT 125.680 130.220 125.910 130.415 ;
        RECT 126.840 130.400 127.170 130.415 ;
        RECT 125.580 129.590 125.910 130.220 ;
        RECT 127.340 130.210 127.570 130.810 ;
        RECT 127.240 129.580 127.570 130.210 ;
        RECT 126.410 128.675 128.490 128.995 ;
        RECT 126.410 128.595 127.480 128.675 ;
        RECT 127.970 128.595 128.490 128.675 ;
        RECT 126.410 128.420 126.650 128.595 ;
        RECT 126.405 128.070 126.655 128.420 ;
        RECT 126.835 127.900 127.475 127.970 ;
        RECT 126.065 127.730 127.475 127.900 ;
        RECT 126.065 127.550 126.235 127.730 ;
        RECT 126.835 127.640 127.475 127.730 ;
        RECT 125.280 127.220 126.235 127.550 ;
        RECT 126.405 127.210 126.655 127.560 ;
        RECT 126.410 127.035 126.650 127.210 ;
        RECT 126.400 126.575 126.650 127.035 ;
        RECT 125.295 126.345 127.505 126.575 ;
        RECT 125.295 126.245 126.275 126.345 ;
        RECT 126.875 126.245 127.505 126.345 ;
        RECT 23.060 121.860 23.560 122.030 ;
        RECT 23.850 121.860 24.350 122.030 ;
        RECT 24.640 121.860 25.140 122.030 ;
        RECT 25.430 121.860 25.930 122.030 ;
        RECT 26.220 121.860 26.720 122.030 ;
        RECT 27.010 121.860 27.510 122.030 ;
        RECT 27.800 121.860 28.300 122.030 ;
        RECT 28.590 121.860 29.090 122.030 ;
        RECT 29.380 121.860 29.880 122.030 ;
        RECT 30.170 121.860 30.670 122.030 ;
        RECT 30.960 121.860 31.460 122.030 ;
        RECT 31.750 121.860 32.250 122.030 ;
        RECT 32.540 121.860 33.040 122.030 ;
        RECT 33.330 121.860 33.830 122.030 ;
        RECT 34.120 121.860 34.620 122.030 ;
        RECT 34.910 121.860 35.410 122.030 ;
        RECT 35.700 121.860 36.200 122.030 ;
        RECT 36.490 121.860 36.990 122.030 ;
        RECT 106.080 121.860 106.580 122.030 ;
        RECT 106.870 121.860 107.370 122.030 ;
        RECT 107.660 121.860 108.160 122.030 ;
        RECT 108.450 121.860 108.950 122.030 ;
        RECT 109.240 121.860 109.740 122.030 ;
        RECT 110.030 121.860 110.530 122.030 ;
        RECT 110.820 121.860 111.320 122.030 ;
        RECT 111.610 121.860 112.110 122.030 ;
        RECT 112.400 121.860 112.900 122.030 ;
        RECT 113.190 121.860 113.690 122.030 ;
        RECT 113.980 121.860 114.480 122.030 ;
        RECT 114.770 121.860 115.270 122.030 ;
        RECT 115.560 121.860 116.060 122.030 ;
        RECT 116.350 121.860 116.850 122.030 ;
        RECT 117.140 121.860 117.640 122.030 ;
        RECT 117.930 121.860 118.430 122.030 ;
        RECT 118.720 121.860 119.220 122.030 ;
        RECT 119.510 121.860 120.010 122.030 ;
        RECT 23.565 117.065 24.065 117.235 ;
        RECT 24.355 117.065 24.855 117.235 ;
        RECT 25.145 117.065 25.645 117.235 ;
        RECT 25.935 117.065 26.435 117.235 ;
        RECT 26.725 117.065 27.225 117.235 ;
        RECT 27.515 117.065 28.015 117.235 ;
        RECT 28.305 117.065 28.805 117.235 ;
        RECT 29.095 117.065 29.595 117.235 ;
        RECT 29.885 117.065 30.385 117.235 ;
        RECT 30.675 117.065 31.175 117.235 ;
        RECT 31.465 117.065 31.965 117.235 ;
        RECT 32.255 117.065 32.755 117.235 ;
        RECT 33.045 117.065 33.545 117.235 ;
        RECT 33.835 117.065 34.335 117.235 ;
        RECT 34.625 117.065 35.125 117.235 ;
        RECT 35.415 117.065 35.915 117.235 ;
        RECT 36.205 117.065 36.705 117.235 ;
        RECT 36.995 117.065 37.495 117.235 ;
        RECT 23.335 106.810 23.505 116.850 ;
        RECT 24.915 106.810 25.085 116.850 ;
        RECT 26.495 106.810 26.665 116.850 ;
        RECT 28.075 106.810 28.245 116.850 ;
        RECT 29.655 106.810 29.825 116.850 ;
        RECT 31.235 106.810 31.405 116.850 ;
        RECT 32.815 106.810 32.985 116.850 ;
        RECT 34.395 106.810 34.565 116.850 ;
        RECT 35.975 106.810 36.145 116.850 ;
        RECT 37.555 106.810 37.725 116.850 ;
        RECT 106.235 116.395 106.735 116.565 ;
        RECT 107.025 116.395 107.525 116.565 ;
        RECT 107.815 116.395 108.315 116.565 ;
        RECT 108.605 116.395 109.105 116.565 ;
        RECT 109.395 116.395 109.895 116.565 ;
        RECT 110.185 116.395 110.685 116.565 ;
        RECT 110.975 116.395 111.475 116.565 ;
        RECT 111.765 116.395 112.265 116.565 ;
        RECT 112.555 116.395 113.055 116.565 ;
        RECT 113.345 116.395 113.845 116.565 ;
        RECT 114.135 116.395 114.635 116.565 ;
        RECT 114.925 116.395 115.425 116.565 ;
        RECT 115.715 116.395 116.215 116.565 ;
        RECT 116.505 116.395 117.005 116.565 ;
        RECT 117.295 116.395 117.795 116.565 ;
        RECT 118.085 116.395 118.585 116.565 ;
        RECT 118.875 116.395 119.375 116.565 ;
        RECT 119.665 116.395 120.165 116.565 ;
        RECT 23.565 106.425 24.065 106.595 ;
        RECT 24.355 106.425 24.855 106.595 ;
        RECT 25.145 106.425 25.645 106.595 ;
        RECT 25.935 106.425 26.435 106.595 ;
        RECT 26.725 106.425 27.225 106.595 ;
        RECT 27.515 106.425 28.015 106.595 ;
        RECT 28.305 106.425 28.805 106.595 ;
        RECT 29.095 106.425 29.595 106.595 ;
        RECT 29.885 106.425 30.385 106.595 ;
        RECT 30.675 106.425 31.175 106.595 ;
        RECT 31.465 106.425 31.965 106.595 ;
        RECT 32.255 106.425 32.755 106.595 ;
        RECT 33.045 106.425 33.545 106.595 ;
        RECT 33.835 106.425 34.335 106.595 ;
        RECT 34.625 106.425 35.125 106.595 ;
        RECT 35.415 106.425 35.915 106.595 ;
        RECT 36.205 106.425 36.705 106.595 ;
        RECT 36.995 106.425 37.495 106.595 ;
        RECT 106.005 106.140 106.175 116.180 ;
        RECT 107.585 106.140 107.755 116.180 ;
        RECT 109.165 106.140 109.335 116.180 ;
        RECT 110.745 106.140 110.915 116.180 ;
        RECT 112.325 106.140 112.495 116.180 ;
        RECT 113.905 106.140 114.075 116.180 ;
        RECT 115.485 106.140 115.655 116.180 ;
        RECT 117.065 106.140 117.235 116.180 ;
        RECT 118.645 106.140 118.815 116.180 ;
        RECT 120.225 106.140 120.395 116.180 ;
        RECT 106.235 105.755 106.735 105.925 ;
        RECT 107.025 105.755 107.525 105.925 ;
        RECT 107.815 105.755 108.315 105.925 ;
        RECT 108.605 105.755 109.105 105.925 ;
        RECT 109.395 105.755 109.895 105.925 ;
        RECT 110.185 105.755 110.685 105.925 ;
        RECT 110.975 105.755 111.475 105.925 ;
        RECT 111.765 105.755 112.265 105.925 ;
        RECT 112.555 105.755 113.055 105.925 ;
        RECT 113.345 105.755 113.845 105.925 ;
        RECT 114.135 105.755 114.635 105.925 ;
        RECT 114.925 105.755 115.425 105.925 ;
        RECT 115.715 105.755 116.215 105.925 ;
        RECT 116.505 105.755 117.005 105.925 ;
        RECT 117.295 105.755 117.795 105.925 ;
        RECT 118.085 105.755 118.585 105.925 ;
        RECT 118.875 105.755 119.375 105.925 ;
        RECT 119.665 105.755 120.165 105.925 ;
        RECT 38.205 104.295 38.795 104.465 ;
        RECT 23.415 103.495 23.915 103.665 ;
        RECT 24.205 103.495 24.705 103.665 ;
        RECT 24.995 103.495 25.495 103.665 ;
        RECT 25.785 103.495 26.285 103.665 ;
        RECT 26.575 103.495 27.075 103.665 ;
        RECT 27.365 103.495 27.865 103.665 ;
        RECT 28.155 103.495 28.655 103.665 ;
        RECT 28.945 103.495 29.445 103.665 ;
        RECT 29.735 103.495 30.235 103.665 ;
        RECT 30.525 103.495 31.025 103.665 ;
        RECT 31.315 103.495 31.815 103.665 ;
        RECT 32.105 103.495 32.605 103.665 ;
        RECT 23.185 98.285 23.355 103.325 ;
        RECT 24.765 98.285 24.935 103.325 ;
        RECT 26.345 98.285 26.515 103.325 ;
        RECT 27.925 98.285 28.095 103.325 ;
        RECT 29.505 98.285 29.675 103.325 ;
        RECT 31.085 98.285 31.255 103.325 ;
        RECT 32.665 98.285 32.835 103.325 ;
        RECT 36.505 102.555 36.675 104.145 ;
        RECT 38.715 103.475 39.045 104.065 ;
        RECT 104.935 103.625 105.525 103.795 ;
        RECT 36.845 103.225 39.045 103.475 ;
        RECT 38.715 102.635 39.045 103.225 ;
        RECT 104.685 102.805 105.015 103.395 ;
        RECT 104.685 102.555 106.885 102.805 ;
        RECT 38.155 102.185 38.765 102.355 ;
        RECT 104.685 101.965 105.015 102.555 ;
        RECT 107.055 101.885 107.225 103.475 ;
        RECT 111.125 102.825 111.625 102.995 ;
        RECT 111.915 102.825 112.415 102.995 ;
        RECT 112.705 102.825 113.205 102.995 ;
        RECT 113.495 102.825 113.995 102.995 ;
        RECT 114.285 102.825 114.785 102.995 ;
        RECT 115.075 102.825 115.575 102.995 ;
        RECT 115.865 102.825 116.365 102.995 ;
        RECT 116.655 102.825 117.155 102.995 ;
        RECT 117.445 102.825 117.945 102.995 ;
        RECT 118.235 102.825 118.735 102.995 ;
        RECT 119.025 102.825 119.525 102.995 ;
        RECT 119.815 102.825 120.315 102.995 ;
        RECT 38.205 101.555 38.815 101.725 ;
        RECT 104.965 101.515 105.575 101.685 ;
        RECT 36.505 99.765 36.675 101.355 ;
        RECT 38.715 100.685 39.045 101.275 ;
        RECT 104.915 100.885 105.525 101.055 ;
        RECT 36.845 100.435 39.045 100.685 ;
        RECT 38.715 99.845 39.045 100.435 ;
        RECT 104.685 100.015 105.015 100.605 ;
        RECT 104.685 99.765 106.885 100.015 ;
        RECT 38.205 99.445 38.795 99.615 ;
        RECT 104.685 99.175 105.015 99.765 ;
        RECT 107.055 99.095 107.225 100.685 ;
        RECT 104.935 98.775 105.525 98.945 ;
        RECT 37.345 98.175 37.685 98.345 ;
        RECT 38.405 98.175 39.325 98.345 ;
        RECT 23.415 97.945 23.915 98.115 ;
        RECT 24.205 97.945 24.705 98.115 ;
        RECT 24.995 97.945 25.495 98.115 ;
        RECT 25.785 97.945 26.285 98.115 ;
        RECT 26.575 97.945 27.075 98.115 ;
        RECT 27.365 97.945 27.865 98.115 ;
        RECT 28.155 97.945 28.655 98.115 ;
        RECT 28.945 97.945 29.445 98.115 ;
        RECT 29.735 97.945 30.235 98.115 ;
        RECT 30.525 97.945 31.025 98.115 ;
        RECT 31.315 97.945 31.815 98.115 ;
        RECT 32.105 97.945 32.605 98.115 ;
        RECT 37.955 97.745 38.125 98.115 ;
        RECT 104.405 97.505 105.325 97.675 ;
        RECT 106.045 97.505 106.385 97.675 ;
        RECT 110.895 97.615 111.065 102.655 ;
        RECT 112.475 97.615 112.645 102.655 ;
        RECT 114.055 97.615 114.225 102.655 ;
        RECT 115.635 97.615 115.805 102.655 ;
        RECT 117.215 97.615 117.385 102.655 ;
        RECT 118.795 97.615 118.965 102.655 ;
        RECT 120.375 97.615 120.545 102.655 ;
        RECT 105.605 97.075 105.775 97.445 ;
        RECT 111.125 97.275 111.625 97.445 ;
        RECT 111.915 97.275 112.415 97.445 ;
        RECT 112.705 97.275 113.205 97.445 ;
        RECT 113.495 97.275 113.995 97.445 ;
        RECT 114.285 97.275 114.785 97.445 ;
        RECT 115.075 97.275 115.575 97.445 ;
        RECT 115.865 97.275 116.365 97.445 ;
        RECT 116.655 97.275 117.155 97.445 ;
        RECT 117.445 97.275 117.945 97.445 ;
        RECT 118.235 97.275 118.735 97.445 ;
        RECT 119.025 97.275 119.525 97.445 ;
        RECT 119.815 97.275 120.315 97.445 ;
        RECT 23.090 92.750 23.260 93.120 ;
        RECT 28.610 92.750 29.110 92.920 ;
        RECT 29.400 92.750 29.900 92.920 ;
        RECT 30.190 92.750 30.690 92.920 ;
        RECT 30.980 92.750 31.480 92.920 ;
        RECT 31.770 92.750 32.270 92.920 ;
        RECT 32.560 92.750 33.060 92.920 ;
        RECT 33.350 92.750 33.850 92.920 ;
        RECT 34.140 92.750 34.640 92.920 ;
        RECT 34.930 92.750 35.430 92.920 ;
        RECT 35.720 92.750 36.220 92.920 ;
        RECT 36.510 92.750 37.010 92.920 ;
        RECT 37.300 92.750 37.800 92.920 ;
        RECT 21.890 92.520 22.810 92.690 ;
        RECT 23.530 92.520 23.870 92.690 ;
        RECT 22.420 91.250 23.010 91.420 ;
        RECT 22.170 90.430 22.500 91.020 ;
        RECT 22.170 90.180 24.370 90.430 ;
        RECT 22.170 89.590 22.500 90.180 ;
        RECT 24.540 89.510 24.710 91.100 ;
        RECT 16.325 89.440 16.965 89.510 ;
        RECT 16.325 89.270 17.735 89.440 ;
        RECT 16.325 89.180 16.965 89.270 ;
        RECT 17.145 88.750 17.395 89.100 ;
        RECT 17.565 89.090 17.735 89.270 ;
        RECT 17.565 88.760 18.520 89.090 ;
        RECT 14.440 88.645 14.780 88.745 ;
        RECT 14.960 88.645 15.480 88.655 ;
        RECT 14.440 88.555 15.480 88.645 ;
        RECT 17.150 88.555 17.390 88.750 ;
        RECT 14.440 88.475 15.830 88.555 ;
        RECT 16.330 88.475 17.390 88.555 ;
        RECT 14.440 88.225 17.390 88.475 ;
        RECT 17.860 88.565 18.400 88.760 ;
        RECT 19.140 88.715 19.880 89.215 ;
        RECT 22.400 89.140 23.010 89.310 ;
        RECT 17.860 88.505 18.510 88.565 ;
        RECT 17.860 88.495 18.520 88.505 ;
        RECT 17.860 88.485 18.970 88.495 ;
        RECT 19.140 88.485 19.890 88.715 ;
        RECT 22.450 88.510 23.060 88.680 ;
        RECT 17.860 88.265 19.890 88.485 ;
        RECT 18.150 88.235 19.890 88.265 ;
        RECT 14.440 88.215 15.480 88.225 ;
        RECT 14.440 88.205 15.010 88.215 ;
        RECT 14.440 88.085 14.780 88.205 ;
        RECT 19.010 88.175 19.890 88.235 ;
        RECT 16.000 86.815 16.330 87.670 ;
        RECT 14.480 86.690 16.330 86.815 ;
        RECT 17.720 86.690 18.050 87.670 ;
        RECT 14.480 86.090 16.230 86.690 ;
        RECT 16.400 86.505 16.730 86.520 ;
        RECT 17.720 86.505 17.950 86.690 ;
        RECT 19.010 86.525 19.600 88.175 ;
        RECT 22.170 87.640 22.500 88.230 ;
        RECT 22.170 87.390 24.370 87.640 ;
        RECT 22.170 86.800 22.500 87.390 ;
        RECT 24.540 86.720 24.710 88.310 ;
        RECT 28.380 87.540 28.550 92.580 ;
        RECT 29.960 87.540 30.130 92.580 ;
        RECT 31.540 87.540 31.710 92.580 ;
        RECT 33.120 87.540 33.290 92.580 ;
        RECT 34.700 87.540 34.870 92.580 ;
        RECT 36.280 87.540 36.450 92.580 ;
        RECT 37.860 87.540 38.030 92.580 ;
        RECT 105.930 92.080 106.430 92.250 ;
        RECT 106.720 92.080 107.220 92.250 ;
        RECT 107.510 92.080 108.010 92.250 ;
        RECT 108.300 92.080 108.800 92.250 ;
        RECT 109.090 92.080 109.590 92.250 ;
        RECT 109.880 92.080 110.380 92.250 ;
        RECT 110.670 92.080 111.170 92.250 ;
        RECT 111.460 92.080 111.960 92.250 ;
        RECT 112.250 92.080 112.750 92.250 ;
        RECT 113.040 92.080 113.540 92.250 ;
        RECT 113.830 92.080 114.330 92.250 ;
        RECT 114.620 92.080 115.120 92.250 ;
        RECT 120.470 92.080 120.640 92.450 ;
        RECT 28.610 87.200 29.110 87.370 ;
        RECT 29.400 87.200 29.900 87.370 ;
        RECT 30.190 87.200 30.690 87.370 ;
        RECT 30.980 87.200 31.480 87.370 ;
        RECT 31.770 87.200 32.270 87.370 ;
        RECT 32.560 87.200 33.060 87.370 ;
        RECT 33.350 87.200 33.850 87.370 ;
        RECT 34.140 87.200 34.640 87.370 ;
        RECT 34.930 87.200 35.430 87.370 ;
        RECT 35.720 87.200 36.220 87.370 ;
        RECT 36.510 87.200 37.010 87.370 ;
        RECT 37.300 87.200 37.800 87.370 ;
        RECT 105.700 86.870 105.870 91.910 ;
        RECT 107.280 86.870 107.450 91.910 ;
        RECT 108.860 86.870 109.030 91.910 ;
        RECT 110.440 86.870 110.610 91.910 ;
        RECT 112.020 86.870 112.190 91.910 ;
        RECT 113.600 86.870 113.770 91.910 ;
        RECT 115.180 86.870 115.350 91.910 ;
        RECT 119.860 91.850 120.200 92.020 ;
        RECT 120.920 91.850 121.840 92.020 ;
        RECT 120.720 90.580 121.310 90.750 ;
        RECT 119.020 88.840 119.190 90.430 ;
        RECT 121.230 89.760 121.560 90.350 ;
        RECT 119.360 89.510 121.560 89.760 ;
        RECT 121.230 88.920 121.560 89.510 ;
        RECT 126.765 88.770 127.405 88.840 ;
        RECT 120.720 88.470 121.330 88.640 ;
        RECT 125.995 88.600 127.405 88.770 ;
        RECT 123.850 88.045 124.590 88.545 ;
        RECT 125.995 88.420 126.165 88.600 ;
        RECT 126.765 88.510 127.405 88.600 ;
        RECT 125.210 88.090 126.165 88.420 ;
        RECT 120.670 87.840 121.280 88.010 ;
        RECT 123.840 87.815 124.590 88.045 ;
        RECT 125.330 87.895 125.870 88.090 ;
        RECT 126.335 88.080 126.585 88.430 ;
        RECT 125.220 87.835 125.870 87.895 ;
        RECT 125.210 87.825 125.870 87.835 ;
        RECT 124.760 87.815 125.870 87.825 ;
        RECT 18.240 86.520 19.600 86.525 ;
        RECT 16.400 86.285 17.950 86.505 ;
        RECT 16.400 86.280 16.730 86.285 ;
        RECT 17.720 86.090 17.950 86.285 ;
        RECT 18.120 86.285 19.600 86.520 ;
        RECT 22.420 86.400 23.010 86.570 ;
        RECT 105.930 86.530 106.430 86.700 ;
        RECT 106.720 86.530 107.220 86.700 ;
        RECT 107.510 86.530 108.010 86.700 ;
        RECT 108.300 86.530 108.800 86.700 ;
        RECT 109.090 86.530 109.590 86.700 ;
        RECT 109.880 86.530 110.380 86.700 ;
        RECT 110.670 86.530 111.170 86.700 ;
        RECT 111.460 86.530 111.960 86.700 ;
        RECT 112.250 86.530 112.750 86.700 ;
        RECT 113.040 86.530 113.540 86.700 ;
        RECT 113.830 86.530 114.330 86.700 ;
        RECT 114.620 86.530 115.120 86.700 ;
        RECT 18.120 86.280 18.450 86.285 ;
        RECT 14.480 86.025 16.330 86.090 ;
        RECT 16.000 85.460 16.330 86.025 ;
        RECT 17.720 85.460 18.050 86.090 ;
        RECT 119.020 86.050 119.190 87.640 ;
        RECT 123.840 87.595 125.870 87.815 ;
        RECT 126.340 87.885 126.580 88.080 ;
        RECT 128.250 87.975 128.770 87.985 ;
        RECT 128.950 87.975 129.290 88.075 ;
        RECT 128.250 87.885 129.290 87.975 ;
        RECT 126.340 87.805 127.400 87.885 ;
        RECT 127.900 87.805 129.290 87.885 ;
        RECT 123.840 87.565 125.580 87.595 ;
        RECT 121.230 86.970 121.560 87.560 ;
        RECT 123.840 87.505 124.720 87.565 ;
        RECT 126.340 87.555 129.290 87.805 ;
        RECT 128.250 87.545 129.290 87.555 ;
        RECT 128.720 87.535 129.290 87.545 ;
        RECT 119.360 86.720 121.560 86.970 ;
        RECT 121.230 86.130 121.560 86.720 ;
        RECT 120.720 85.730 121.310 85.900 ;
        RECT 124.130 85.855 124.720 87.505 ;
        RECT 128.950 87.415 129.290 87.535 ;
        RECT 125.680 86.020 126.010 87.000 ;
        RECT 127.400 86.145 127.730 87.000 ;
        RECT 127.400 86.020 129.250 86.145 ;
        RECT 124.130 85.850 125.490 85.855 ;
        RECT 124.130 85.615 125.610 85.850 ;
        RECT 125.280 85.610 125.610 85.615 ;
        RECT 125.780 85.835 126.010 86.020 ;
        RECT 127.000 85.835 127.330 85.850 ;
        RECT 125.780 85.615 127.330 85.835 ;
        RECT 125.780 85.420 126.010 85.615 ;
        RECT 127.000 85.610 127.330 85.615 ;
        RECT 127.500 85.420 129.250 86.020 ;
        RECT 125.680 84.790 126.010 85.420 ;
        RECT 127.400 85.355 129.250 85.420 ;
        RECT 127.400 84.790 127.730 85.355 ;
        RECT 23.720 84.270 24.220 84.440 ;
        RECT 24.510 84.270 25.010 84.440 ;
        RECT 25.300 84.270 25.800 84.440 ;
        RECT 26.090 84.270 26.590 84.440 ;
        RECT 26.880 84.270 27.380 84.440 ;
        RECT 27.670 84.270 28.170 84.440 ;
        RECT 28.460 84.270 28.960 84.440 ;
        RECT 29.250 84.270 29.750 84.440 ;
        RECT 30.040 84.270 30.540 84.440 ;
        RECT 30.830 84.270 31.330 84.440 ;
        RECT 31.620 84.270 32.120 84.440 ;
        RECT 32.410 84.270 32.910 84.440 ;
        RECT 33.200 84.270 33.700 84.440 ;
        RECT 33.990 84.270 34.490 84.440 ;
        RECT 34.780 84.270 35.280 84.440 ;
        RECT 35.570 84.270 36.070 84.440 ;
        RECT 36.360 84.270 36.860 84.440 ;
        RECT 37.150 84.270 37.650 84.440 ;
        RECT 16.160 83.335 16.490 83.560 ;
        RECT 15.780 82.775 16.490 83.335 ;
        RECT 16.160 82.580 16.490 82.775 ;
        RECT 17.820 82.590 18.150 83.570 ;
        RECT 16.160 81.980 16.390 82.580 ;
        RECT 16.560 82.375 16.890 82.410 ;
        RECT 17.820 82.375 18.050 82.590 ;
        RECT 16.560 82.185 18.050 82.375 ;
        RECT 16.560 82.170 16.890 82.185 ;
        RECT 17.820 81.990 18.050 82.185 ;
        RECT 18.220 82.415 18.550 82.420 ;
        RECT 18.860 82.415 19.690 82.505 ;
        RECT 18.220 82.185 19.690 82.415 ;
        RECT 18.220 82.180 18.550 82.185 ;
        RECT 16.160 81.350 16.490 81.980 ;
        RECT 17.820 81.360 18.150 81.990 ;
        RECT 18.860 81.985 19.690 82.185 ;
        RECT 15.240 80.445 17.320 80.765 ;
        RECT 15.240 80.365 15.760 80.445 ;
        RECT 16.250 80.365 17.320 80.445 ;
        RECT 17.080 80.190 17.320 80.365 ;
        RECT 17.075 79.840 17.325 80.190 ;
        RECT 16.255 79.670 16.895 79.740 ;
        RECT 16.255 79.500 17.665 79.670 ;
        RECT 16.255 79.410 16.895 79.500 ;
        RECT 17.075 78.980 17.325 79.330 ;
        RECT 17.495 79.320 17.665 79.500 ;
        RECT 17.495 78.990 18.450 79.320 ;
        RECT 17.080 78.805 17.320 78.980 ;
        RECT 17.080 78.345 17.330 78.805 ;
        RECT 16.225 78.115 18.435 78.345 ;
        RECT 16.225 78.015 16.855 78.115 ;
        RECT 17.455 78.015 18.435 78.115 ;
        RECT 23.490 74.015 23.660 84.055 ;
        RECT 25.070 74.015 25.240 84.055 ;
        RECT 26.650 74.015 26.820 84.055 ;
        RECT 28.230 74.015 28.400 84.055 ;
        RECT 29.810 74.015 29.980 84.055 ;
        RECT 31.390 74.015 31.560 84.055 ;
        RECT 32.970 74.015 33.140 84.055 ;
        RECT 34.550 74.015 34.720 84.055 ;
        RECT 36.130 74.015 36.300 84.055 ;
        RECT 37.710 74.015 37.880 84.055 ;
        RECT 106.080 83.600 106.580 83.770 ;
        RECT 106.870 83.600 107.370 83.770 ;
        RECT 107.660 83.600 108.160 83.770 ;
        RECT 108.450 83.600 108.950 83.770 ;
        RECT 109.240 83.600 109.740 83.770 ;
        RECT 110.030 83.600 110.530 83.770 ;
        RECT 110.820 83.600 111.320 83.770 ;
        RECT 111.610 83.600 112.110 83.770 ;
        RECT 112.400 83.600 112.900 83.770 ;
        RECT 113.190 83.600 113.690 83.770 ;
        RECT 113.980 83.600 114.480 83.770 ;
        RECT 114.770 83.600 115.270 83.770 ;
        RECT 115.560 83.600 116.060 83.770 ;
        RECT 116.350 83.600 116.850 83.770 ;
        RECT 117.140 83.600 117.640 83.770 ;
        RECT 117.930 83.600 118.430 83.770 ;
        RECT 118.720 83.600 119.220 83.770 ;
        RECT 119.510 83.600 120.010 83.770 ;
        RECT 23.720 73.630 24.220 73.800 ;
        RECT 24.510 73.630 25.010 73.800 ;
        RECT 25.300 73.630 25.800 73.800 ;
        RECT 26.090 73.630 26.590 73.800 ;
        RECT 26.880 73.630 27.380 73.800 ;
        RECT 27.670 73.630 28.170 73.800 ;
        RECT 28.460 73.630 28.960 73.800 ;
        RECT 29.250 73.630 29.750 73.800 ;
        RECT 30.040 73.630 30.540 73.800 ;
        RECT 30.830 73.630 31.330 73.800 ;
        RECT 31.620 73.630 32.120 73.800 ;
        RECT 32.410 73.630 32.910 73.800 ;
        RECT 33.200 73.630 33.700 73.800 ;
        RECT 33.990 73.630 34.490 73.800 ;
        RECT 34.780 73.630 35.280 73.800 ;
        RECT 35.570 73.630 36.070 73.800 ;
        RECT 36.360 73.630 36.860 73.800 ;
        RECT 37.150 73.630 37.650 73.800 ;
        RECT 105.850 73.345 106.020 83.385 ;
        RECT 107.430 73.345 107.600 83.385 ;
        RECT 109.010 73.345 109.180 83.385 ;
        RECT 110.590 73.345 110.760 83.385 ;
        RECT 112.170 73.345 112.340 83.385 ;
        RECT 113.750 73.345 113.920 83.385 ;
        RECT 115.330 73.345 115.500 83.385 ;
        RECT 116.910 73.345 117.080 83.385 ;
        RECT 118.490 73.345 118.660 83.385 ;
        RECT 120.070 73.345 120.240 83.385 ;
        RECT 125.580 81.920 125.910 82.900 ;
        RECT 124.040 81.745 124.870 81.835 ;
        RECT 125.180 81.745 125.510 81.750 ;
        RECT 124.040 81.515 125.510 81.745 ;
        RECT 124.040 81.315 124.870 81.515 ;
        RECT 125.180 81.510 125.510 81.515 ;
        RECT 125.680 81.705 125.910 81.920 ;
        RECT 127.240 82.665 127.570 82.890 ;
        RECT 127.240 82.105 127.950 82.665 ;
        RECT 127.240 81.910 127.570 82.105 ;
        RECT 126.840 81.705 127.170 81.740 ;
        RECT 125.680 81.515 127.170 81.705 ;
        RECT 125.680 81.320 125.910 81.515 ;
        RECT 126.840 81.500 127.170 81.515 ;
        RECT 125.580 80.690 125.910 81.320 ;
        RECT 127.340 81.310 127.570 81.910 ;
        RECT 127.240 80.680 127.570 81.310 ;
        RECT 126.410 79.775 128.490 80.095 ;
        RECT 126.410 79.695 127.480 79.775 ;
        RECT 127.970 79.695 128.490 79.775 ;
        RECT 126.410 79.520 126.650 79.695 ;
        RECT 126.405 79.170 126.655 79.520 ;
        RECT 126.835 79.000 127.475 79.070 ;
        RECT 126.065 78.830 127.475 79.000 ;
        RECT 126.065 78.650 126.235 78.830 ;
        RECT 126.835 78.740 127.475 78.830 ;
        RECT 125.280 78.320 126.235 78.650 ;
        RECT 126.405 78.310 126.655 78.660 ;
        RECT 126.410 78.135 126.650 78.310 ;
        RECT 126.400 77.675 126.650 78.135 ;
        RECT 125.295 77.445 127.505 77.675 ;
        RECT 125.295 77.345 126.275 77.445 ;
        RECT 126.875 77.345 127.505 77.445 ;
        RECT 106.080 72.960 106.580 73.130 ;
        RECT 106.870 72.960 107.370 73.130 ;
        RECT 107.660 72.960 108.160 73.130 ;
        RECT 108.450 72.960 108.950 73.130 ;
        RECT 109.240 72.960 109.740 73.130 ;
        RECT 110.030 72.960 110.530 73.130 ;
        RECT 110.820 72.960 111.320 73.130 ;
        RECT 111.610 72.960 112.110 73.130 ;
        RECT 112.400 72.960 112.900 73.130 ;
        RECT 113.190 72.960 113.690 73.130 ;
        RECT 113.980 72.960 114.480 73.130 ;
        RECT 114.770 72.960 115.270 73.130 ;
        RECT 115.560 72.960 116.060 73.130 ;
        RECT 116.350 72.960 116.850 73.130 ;
        RECT 117.140 72.960 117.640 73.130 ;
        RECT 117.930 72.960 118.430 73.130 ;
        RECT 118.720 72.960 119.220 73.130 ;
        RECT 119.510 72.960 120.010 73.130 ;
        RECT 23.235 66.495 23.735 66.665 ;
        RECT 24.025 66.495 24.525 66.665 ;
        RECT 24.815 66.495 25.315 66.665 ;
        RECT 25.605 66.495 26.105 66.665 ;
        RECT 26.395 66.495 26.895 66.665 ;
        RECT 27.185 66.495 27.685 66.665 ;
        RECT 27.975 66.495 28.475 66.665 ;
        RECT 28.765 66.495 29.265 66.665 ;
        RECT 29.555 66.495 30.055 66.665 ;
        RECT 30.345 66.495 30.845 66.665 ;
        RECT 31.135 66.495 31.635 66.665 ;
        RECT 31.925 66.495 32.425 66.665 ;
        RECT 32.715 66.495 33.215 66.665 ;
        RECT 33.505 66.495 34.005 66.665 ;
        RECT 34.295 66.495 34.795 66.665 ;
        RECT 35.085 66.495 35.585 66.665 ;
        RECT 35.875 66.495 36.375 66.665 ;
        RECT 36.665 66.495 37.165 66.665 ;
        RECT 105.575 66.495 106.075 66.665 ;
        RECT 106.365 66.495 106.865 66.665 ;
        RECT 107.155 66.495 107.655 66.665 ;
        RECT 107.945 66.495 108.445 66.665 ;
        RECT 108.735 66.495 109.235 66.665 ;
        RECT 109.525 66.495 110.025 66.665 ;
        RECT 110.315 66.495 110.815 66.665 ;
        RECT 111.105 66.495 111.605 66.665 ;
        RECT 111.895 66.495 112.395 66.665 ;
        RECT 112.685 66.495 113.185 66.665 ;
        RECT 113.475 66.495 113.975 66.665 ;
        RECT 114.265 66.495 114.765 66.665 ;
        RECT 115.055 66.495 115.555 66.665 ;
        RECT 115.845 66.495 116.345 66.665 ;
        RECT 116.635 66.495 117.135 66.665 ;
        RECT 117.425 66.495 117.925 66.665 ;
        RECT 118.215 66.495 118.715 66.665 ;
        RECT 119.005 66.495 119.505 66.665 ;
        RECT 23.005 56.240 23.175 66.280 ;
        RECT 24.585 56.240 24.755 66.280 ;
        RECT 26.165 56.240 26.335 66.280 ;
        RECT 27.745 56.240 27.915 66.280 ;
        RECT 29.325 56.240 29.495 66.280 ;
        RECT 30.905 56.240 31.075 66.280 ;
        RECT 32.485 56.240 32.655 66.280 ;
        RECT 34.065 56.240 34.235 66.280 ;
        RECT 35.645 56.240 35.815 66.280 ;
        RECT 37.225 56.240 37.395 66.280 ;
        RECT 105.345 56.240 105.515 66.280 ;
        RECT 106.925 56.240 107.095 66.280 ;
        RECT 108.505 56.240 108.675 66.280 ;
        RECT 110.085 56.240 110.255 66.280 ;
        RECT 111.665 56.240 111.835 66.280 ;
        RECT 113.245 56.240 113.415 66.280 ;
        RECT 114.825 56.240 114.995 66.280 ;
        RECT 116.405 56.240 116.575 66.280 ;
        RECT 117.985 56.240 118.155 66.280 ;
        RECT 119.565 56.240 119.735 66.280 ;
        RECT 23.235 55.855 23.735 56.025 ;
        RECT 24.025 55.855 24.525 56.025 ;
        RECT 24.815 55.855 25.315 56.025 ;
        RECT 25.605 55.855 26.105 56.025 ;
        RECT 26.395 55.855 26.895 56.025 ;
        RECT 27.185 55.855 27.685 56.025 ;
        RECT 27.975 55.855 28.475 56.025 ;
        RECT 28.765 55.855 29.265 56.025 ;
        RECT 29.555 55.855 30.055 56.025 ;
        RECT 30.345 55.855 30.845 56.025 ;
        RECT 31.135 55.855 31.635 56.025 ;
        RECT 31.925 55.855 32.425 56.025 ;
        RECT 32.715 55.855 33.215 56.025 ;
        RECT 33.505 55.855 34.005 56.025 ;
        RECT 34.295 55.855 34.795 56.025 ;
        RECT 35.085 55.855 35.585 56.025 ;
        RECT 35.875 55.855 36.375 56.025 ;
        RECT 36.665 55.855 37.165 56.025 ;
        RECT 105.575 55.855 106.075 56.025 ;
        RECT 106.365 55.855 106.865 56.025 ;
        RECT 107.155 55.855 107.655 56.025 ;
        RECT 107.945 55.855 108.445 56.025 ;
        RECT 108.735 55.855 109.235 56.025 ;
        RECT 109.525 55.855 110.025 56.025 ;
        RECT 110.315 55.855 110.815 56.025 ;
        RECT 111.105 55.855 111.605 56.025 ;
        RECT 111.895 55.855 112.395 56.025 ;
        RECT 112.685 55.855 113.185 56.025 ;
        RECT 113.475 55.855 113.975 56.025 ;
        RECT 114.265 55.855 114.765 56.025 ;
        RECT 115.055 55.855 115.555 56.025 ;
        RECT 115.845 55.855 116.345 56.025 ;
        RECT 116.635 55.855 117.135 56.025 ;
        RECT 117.425 55.855 117.925 56.025 ;
        RECT 118.215 55.855 118.715 56.025 ;
        RECT 119.005 55.855 119.505 56.025 ;
        RECT 37.875 53.725 38.465 53.895 ;
        RECT 104.275 53.725 104.865 53.895 ;
        RECT 23.085 52.925 23.585 53.095 ;
        RECT 23.875 52.925 24.375 53.095 ;
        RECT 24.665 52.925 25.165 53.095 ;
        RECT 25.455 52.925 25.955 53.095 ;
        RECT 26.245 52.925 26.745 53.095 ;
        RECT 27.035 52.925 27.535 53.095 ;
        RECT 27.825 52.925 28.325 53.095 ;
        RECT 28.615 52.925 29.115 53.095 ;
        RECT 29.405 52.925 29.905 53.095 ;
        RECT 30.195 52.925 30.695 53.095 ;
        RECT 30.985 52.925 31.485 53.095 ;
        RECT 31.775 52.925 32.275 53.095 ;
        RECT 22.855 47.715 23.025 52.755 ;
        RECT 24.435 47.715 24.605 52.755 ;
        RECT 26.015 47.715 26.185 52.755 ;
        RECT 27.595 47.715 27.765 52.755 ;
        RECT 29.175 47.715 29.345 52.755 ;
        RECT 30.755 47.715 30.925 52.755 ;
        RECT 32.335 47.715 32.505 52.755 ;
        RECT 36.175 51.985 36.345 53.575 ;
        RECT 38.385 52.905 38.715 53.495 ;
        RECT 36.515 52.655 38.715 52.905 ;
        RECT 38.385 52.065 38.715 52.655 ;
        RECT 104.025 52.905 104.355 53.495 ;
        RECT 104.025 52.655 106.225 52.905 ;
        RECT 104.025 52.065 104.355 52.655 ;
        RECT 106.395 51.985 106.565 53.575 ;
        RECT 110.465 52.925 110.965 53.095 ;
        RECT 111.255 52.925 111.755 53.095 ;
        RECT 112.045 52.925 112.545 53.095 ;
        RECT 112.835 52.925 113.335 53.095 ;
        RECT 113.625 52.925 114.125 53.095 ;
        RECT 114.415 52.925 114.915 53.095 ;
        RECT 115.205 52.925 115.705 53.095 ;
        RECT 115.995 52.925 116.495 53.095 ;
        RECT 116.785 52.925 117.285 53.095 ;
        RECT 117.575 52.925 118.075 53.095 ;
        RECT 118.365 52.925 118.865 53.095 ;
        RECT 119.155 52.925 119.655 53.095 ;
        RECT 37.825 51.615 38.435 51.785 ;
        RECT 104.305 51.615 104.915 51.785 ;
        RECT 37.875 50.985 38.485 51.155 ;
        RECT 104.255 50.985 104.865 51.155 ;
        RECT 36.175 49.195 36.345 50.785 ;
        RECT 38.385 50.115 38.715 50.705 ;
        RECT 36.515 49.865 38.715 50.115 ;
        RECT 38.385 49.275 38.715 49.865 ;
        RECT 104.025 50.115 104.355 50.705 ;
        RECT 104.025 49.865 106.225 50.115 ;
        RECT 104.025 49.275 104.355 49.865 ;
        RECT 106.395 49.195 106.565 50.785 ;
        RECT 37.875 48.875 38.465 49.045 ;
        RECT 104.275 48.875 104.865 49.045 ;
        RECT 37.015 47.605 37.355 47.775 ;
        RECT 38.075 47.605 38.995 47.775 ;
        RECT 103.745 47.605 104.665 47.775 ;
        RECT 105.385 47.605 105.725 47.775 ;
        RECT 110.235 47.715 110.405 52.755 ;
        RECT 111.815 47.715 111.985 52.755 ;
        RECT 113.395 47.715 113.565 52.755 ;
        RECT 114.975 47.715 115.145 52.755 ;
        RECT 116.555 47.715 116.725 52.755 ;
        RECT 118.135 47.715 118.305 52.755 ;
        RECT 119.715 47.715 119.885 52.755 ;
        RECT 23.085 47.375 23.585 47.545 ;
        RECT 23.875 47.375 24.375 47.545 ;
        RECT 24.665 47.375 25.165 47.545 ;
        RECT 25.455 47.375 25.955 47.545 ;
        RECT 26.245 47.375 26.745 47.545 ;
        RECT 27.035 47.375 27.535 47.545 ;
        RECT 27.825 47.375 28.325 47.545 ;
        RECT 28.615 47.375 29.115 47.545 ;
        RECT 29.405 47.375 29.905 47.545 ;
        RECT 30.195 47.375 30.695 47.545 ;
        RECT 30.985 47.375 31.485 47.545 ;
        RECT 31.775 47.375 32.275 47.545 ;
        RECT 37.625 47.175 37.795 47.545 ;
        RECT 104.945 47.175 105.115 47.545 ;
        RECT 110.465 47.375 110.965 47.545 ;
        RECT 111.255 47.375 111.755 47.545 ;
        RECT 112.045 47.375 112.545 47.545 ;
        RECT 112.835 47.375 113.335 47.545 ;
        RECT 113.625 47.375 114.125 47.545 ;
        RECT 114.415 47.375 114.915 47.545 ;
        RECT 115.205 47.375 115.705 47.545 ;
        RECT 115.995 47.375 116.495 47.545 ;
        RECT 116.785 47.375 117.285 47.545 ;
        RECT 117.575 47.375 118.075 47.545 ;
        RECT 118.365 47.375 118.865 47.545 ;
        RECT 119.155 47.375 119.655 47.545 ;
        RECT 22.760 42.180 22.930 42.550 ;
        RECT 28.280 42.180 28.780 42.350 ;
        RECT 29.070 42.180 29.570 42.350 ;
        RECT 29.860 42.180 30.360 42.350 ;
        RECT 30.650 42.180 31.150 42.350 ;
        RECT 31.440 42.180 31.940 42.350 ;
        RECT 32.230 42.180 32.730 42.350 ;
        RECT 33.020 42.180 33.520 42.350 ;
        RECT 33.810 42.180 34.310 42.350 ;
        RECT 34.600 42.180 35.100 42.350 ;
        RECT 35.390 42.180 35.890 42.350 ;
        RECT 36.180 42.180 36.680 42.350 ;
        RECT 36.970 42.180 37.470 42.350 ;
        RECT 105.270 42.180 105.770 42.350 ;
        RECT 106.060 42.180 106.560 42.350 ;
        RECT 106.850 42.180 107.350 42.350 ;
        RECT 107.640 42.180 108.140 42.350 ;
        RECT 108.430 42.180 108.930 42.350 ;
        RECT 109.220 42.180 109.720 42.350 ;
        RECT 110.010 42.180 110.510 42.350 ;
        RECT 110.800 42.180 111.300 42.350 ;
        RECT 111.590 42.180 112.090 42.350 ;
        RECT 112.380 42.180 112.880 42.350 ;
        RECT 113.170 42.180 113.670 42.350 ;
        RECT 113.960 42.180 114.460 42.350 ;
        RECT 119.810 42.180 119.980 42.550 ;
        RECT 21.560 41.950 22.480 42.120 ;
        RECT 23.200 41.950 23.540 42.120 ;
        RECT 22.090 40.680 22.680 40.850 ;
        RECT 21.840 39.860 22.170 40.450 ;
        RECT 21.840 39.610 24.040 39.860 ;
        RECT 21.840 39.020 22.170 39.610 ;
        RECT 24.210 38.940 24.380 40.530 ;
        RECT 15.995 38.870 16.635 38.940 ;
        RECT 15.995 38.700 17.405 38.870 ;
        RECT 15.995 38.610 16.635 38.700 ;
        RECT 16.815 38.180 17.065 38.530 ;
        RECT 17.235 38.520 17.405 38.700 ;
        RECT 17.235 38.190 18.190 38.520 ;
        RECT 14.110 38.075 14.450 38.175 ;
        RECT 14.630 38.075 15.150 38.085 ;
        RECT 14.110 37.985 15.150 38.075 ;
        RECT 16.820 37.985 17.060 38.180 ;
        RECT 14.110 37.905 15.500 37.985 ;
        RECT 16.000 37.905 17.060 37.985 ;
        RECT 14.110 37.655 17.060 37.905 ;
        RECT 17.530 37.995 18.070 38.190 ;
        RECT 18.810 38.145 19.550 38.645 ;
        RECT 22.070 38.570 22.680 38.740 ;
        RECT 17.530 37.935 18.180 37.995 ;
        RECT 17.530 37.925 18.190 37.935 ;
        RECT 17.530 37.915 18.640 37.925 ;
        RECT 18.810 37.915 19.560 38.145 ;
        RECT 22.120 37.940 22.730 38.110 ;
        RECT 17.530 37.695 19.560 37.915 ;
        RECT 17.820 37.665 19.560 37.695 ;
        RECT 14.110 37.645 15.150 37.655 ;
        RECT 14.110 37.635 14.680 37.645 ;
        RECT 14.110 37.515 14.450 37.635 ;
        RECT 18.680 37.605 19.560 37.665 ;
        RECT 15.670 36.245 16.000 37.100 ;
        RECT 14.150 36.120 16.000 36.245 ;
        RECT 17.390 36.120 17.720 37.100 ;
        RECT 14.150 35.520 15.900 36.120 ;
        RECT 16.070 35.935 16.400 35.950 ;
        RECT 17.390 35.935 17.620 36.120 ;
        RECT 18.680 35.955 19.270 37.605 ;
        RECT 21.840 37.070 22.170 37.660 ;
        RECT 21.840 36.820 24.040 37.070 ;
        RECT 21.840 36.230 22.170 36.820 ;
        RECT 24.210 36.150 24.380 37.740 ;
        RECT 28.050 36.970 28.220 42.010 ;
        RECT 29.630 36.970 29.800 42.010 ;
        RECT 31.210 36.970 31.380 42.010 ;
        RECT 32.790 36.970 32.960 42.010 ;
        RECT 34.370 36.970 34.540 42.010 ;
        RECT 35.950 36.970 36.120 42.010 ;
        RECT 37.530 36.970 37.700 42.010 ;
        RECT 105.040 36.970 105.210 42.010 ;
        RECT 106.620 36.970 106.790 42.010 ;
        RECT 108.200 36.970 108.370 42.010 ;
        RECT 109.780 36.970 109.950 42.010 ;
        RECT 111.360 36.970 111.530 42.010 ;
        RECT 112.940 36.970 113.110 42.010 ;
        RECT 114.520 36.970 114.690 42.010 ;
        RECT 119.200 41.950 119.540 42.120 ;
        RECT 120.260 41.950 121.180 42.120 ;
        RECT 120.060 40.680 120.650 40.850 ;
        RECT 118.360 38.940 118.530 40.530 ;
        RECT 120.570 39.860 120.900 40.450 ;
        RECT 118.700 39.610 120.900 39.860 ;
        RECT 120.570 39.020 120.900 39.610 ;
        RECT 126.105 38.870 126.745 38.940 ;
        RECT 120.060 38.570 120.670 38.740 ;
        RECT 125.335 38.700 126.745 38.870 ;
        RECT 123.190 38.145 123.930 38.645 ;
        RECT 125.335 38.520 125.505 38.700 ;
        RECT 126.105 38.610 126.745 38.700 ;
        RECT 124.550 38.190 125.505 38.520 ;
        RECT 120.010 37.940 120.620 38.110 ;
        RECT 123.180 37.915 123.930 38.145 ;
        RECT 124.670 37.995 125.210 38.190 ;
        RECT 125.675 38.180 125.925 38.530 ;
        RECT 124.560 37.935 125.210 37.995 ;
        RECT 124.550 37.925 125.210 37.935 ;
        RECT 124.100 37.915 125.210 37.925 ;
        RECT 28.280 36.630 28.780 36.800 ;
        RECT 29.070 36.630 29.570 36.800 ;
        RECT 29.860 36.630 30.360 36.800 ;
        RECT 30.650 36.630 31.150 36.800 ;
        RECT 31.440 36.630 31.940 36.800 ;
        RECT 32.230 36.630 32.730 36.800 ;
        RECT 33.020 36.630 33.520 36.800 ;
        RECT 33.810 36.630 34.310 36.800 ;
        RECT 34.600 36.630 35.100 36.800 ;
        RECT 35.390 36.630 35.890 36.800 ;
        RECT 36.180 36.630 36.680 36.800 ;
        RECT 36.970 36.630 37.470 36.800 ;
        RECT 105.270 36.630 105.770 36.800 ;
        RECT 106.060 36.630 106.560 36.800 ;
        RECT 106.850 36.630 107.350 36.800 ;
        RECT 107.640 36.630 108.140 36.800 ;
        RECT 108.430 36.630 108.930 36.800 ;
        RECT 109.220 36.630 109.720 36.800 ;
        RECT 110.010 36.630 110.510 36.800 ;
        RECT 110.800 36.630 111.300 36.800 ;
        RECT 111.590 36.630 112.090 36.800 ;
        RECT 112.380 36.630 112.880 36.800 ;
        RECT 113.170 36.630 113.670 36.800 ;
        RECT 113.960 36.630 114.460 36.800 ;
        RECT 118.360 36.150 118.530 37.740 ;
        RECT 123.180 37.695 125.210 37.915 ;
        RECT 125.680 37.985 125.920 38.180 ;
        RECT 127.590 38.075 128.110 38.085 ;
        RECT 128.290 38.075 128.630 38.175 ;
        RECT 127.590 37.985 128.630 38.075 ;
        RECT 125.680 37.905 126.740 37.985 ;
        RECT 127.240 37.905 128.630 37.985 ;
        RECT 123.180 37.665 124.920 37.695 ;
        RECT 120.570 37.070 120.900 37.660 ;
        RECT 123.180 37.605 124.060 37.665 ;
        RECT 125.680 37.655 128.630 37.905 ;
        RECT 127.590 37.645 128.630 37.655 ;
        RECT 128.060 37.635 128.630 37.645 ;
        RECT 118.700 36.820 120.900 37.070 ;
        RECT 120.570 36.230 120.900 36.820 ;
        RECT 17.910 35.950 19.270 35.955 ;
        RECT 16.070 35.715 17.620 35.935 ;
        RECT 16.070 35.710 16.400 35.715 ;
        RECT 17.390 35.520 17.620 35.715 ;
        RECT 17.790 35.715 19.270 35.950 ;
        RECT 22.090 35.830 22.680 36.000 ;
        RECT 120.060 35.830 120.650 36.000 ;
        RECT 123.470 35.955 124.060 37.605 ;
        RECT 128.290 37.515 128.630 37.635 ;
        RECT 125.020 36.120 125.350 37.100 ;
        RECT 126.740 36.245 127.070 37.100 ;
        RECT 126.740 36.120 128.590 36.245 ;
        RECT 123.470 35.950 124.830 35.955 ;
        RECT 123.470 35.715 124.950 35.950 ;
        RECT 17.790 35.710 18.120 35.715 ;
        RECT 124.620 35.710 124.950 35.715 ;
        RECT 125.120 35.935 125.350 36.120 ;
        RECT 126.340 35.935 126.670 35.950 ;
        RECT 125.120 35.715 126.670 35.935 ;
        RECT 125.120 35.520 125.350 35.715 ;
        RECT 126.340 35.710 126.670 35.715 ;
        RECT 126.840 35.520 128.590 36.120 ;
        RECT 14.150 35.455 16.000 35.520 ;
        RECT 15.670 34.890 16.000 35.455 ;
        RECT 17.390 34.890 17.720 35.520 ;
        RECT 125.020 34.890 125.350 35.520 ;
        RECT 126.740 35.455 128.590 35.520 ;
        RECT 126.740 34.890 127.070 35.455 ;
        RECT 23.390 33.700 23.890 33.870 ;
        RECT 24.180 33.700 24.680 33.870 ;
        RECT 24.970 33.700 25.470 33.870 ;
        RECT 25.760 33.700 26.260 33.870 ;
        RECT 26.550 33.700 27.050 33.870 ;
        RECT 27.340 33.700 27.840 33.870 ;
        RECT 28.130 33.700 28.630 33.870 ;
        RECT 28.920 33.700 29.420 33.870 ;
        RECT 29.710 33.700 30.210 33.870 ;
        RECT 30.500 33.700 31.000 33.870 ;
        RECT 31.290 33.700 31.790 33.870 ;
        RECT 32.080 33.700 32.580 33.870 ;
        RECT 32.870 33.700 33.370 33.870 ;
        RECT 33.660 33.700 34.160 33.870 ;
        RECT 34.450 33.700 34.950 33.870 ;
        RECT 35.240 33.700 35.740 33.870 ;
        RECT 36.030 33.700 36.530 33.870 ;
        RECT 36.820 33.700 37.320 33.870 ;
        RECT 105.420 33.700 105.920 33.870 ;
        RECT 106.210 33.700 106.710 33.870 ;
        RECT 107.000 33.700 107.500 33.870 ;
        RECT 107.790 33.700 108.290 33.870 ;
        RECT 108.580 33.700 109.080 33.870 ;
        RECT 109.370 33.700 109.870 33.870 ;
        RECT 110.160 33.700 110.660 33.870 ;
        RECT 110.950 33.700 111.450 33.870 ;
        RECT 111.740 33.700 112.240 33.870 ;
        RECT 112.530 33.700 113.030 33.870 ;
        RECT 113.320 33.700 113.820 33.870 ;
        RECT 114.110 33.700 114.610 33.870 ;
        RECT 114.900 33.700 115.400 33.870 ;
        RECT 115.690 33.700 116.190 33.870 ;
        RECT 116.480 33.700 116.980 33.870 ;
        RECT 117.270 33.700 117.770 33.870 ;
        RECT 118.060 33.700 118.560 33.870 ;
        RECT 118.850 33.700 119.350 33.870 ;
        RECT 15.830 32.765 16.160 32.990 ;
        RECT 15.450 32.205 16.160 32.765 ;
        RECT 15.830 32.010 16.160 32.205 ;
        RECT 17.490 32.020 17.820 33.000 ;
        RECT 15.830 31.410 16.060 32.010 ;
        RECT 16.230 31.805 16.560 31.840 ;
        RECT 17.490 31.805 17.720 32.020 ;
        RECT 16.230 31.615 17.720 31.805 ;
        RECT 16.230 31.600 16.560 31.615 ;
        RECT 17.490 31.420 17.720 31.615 ;
        RECT 17.890 31.845 18.220 31.850 ;
        RECT 18.530 31.845 19.360 31.935 ;
        RECT 17.890 31.615 19.360 31.845 ;
        RECT 17.890 31.610 18.220 31.615 ;
        RECT 15.830 30.780 16.160 31.410 ;
        RECT 17.490 30.790 17.820 31.420 ;
        RECT 18.530 31.415 19.360 31.615 ;
        RECT 14.910 29.875 16.990 30.195 ;
        RECT 14.910 29.795 15.430 29.875 ;
        RECT 15.920 29.795 16.990 29.875 ;
        RECT 16.750 29.620 16.990 29.795 ;
        RECT 16.745 29.270 16.995 29.620 ;
        RECT 15.925 29.100 16.565 29.170 ;
        RECT 15.925 28.930 17.335 29.100 ;
        RECT 15.925 28.840 16.565 28.930 ;
        RECT 16.745 28.410 16.995 28.760 ;
        RECT 17.165 28.750 17.335 28.930 ;
        RECT 17.165 28.420 18.120 28.750 ;
        RECT 16.750 28.235 16.990 28.410 ;
        RECT 16.750 27.775 17.000 28.235 ;
        RECT 15.895 27.545 18.105 27.775 ;
        RECT 15.895 27.445 16.525 27.545 ;
        RECT 17.125 27.445 18.105 27.545 ;
        RECT 23.160 23.445 23.330 33.485 ;
        RECT 24.740 23.445 24.910 33.485 ;
        RECT 26.320 23.445 26.490 33.485 ;
        RECT 27.900 23.445 28.070 33.485 ;
        RECT 29.480 23.445 29.650 33.485 ;
        RECT 31.060 23.445 31.230 33.485 ;
        RECT 32.640 23.445 32.810 33.485 ;
        RECT 34.220 23.445 34.390 33.485 ;
        RECT 35.800 23.445 35.970 33.485 ;
        RECT 37.380 23.445 37.550 33.485 ;
        RECT 105.190 23.445 105.360 33.485 ;
        RECT 106.770 23.445 106.940 33.485 ;
        RECT 108.350 23.445 108.520 33.485 ;
        RECT 109.930 23.445 110.100 33.485 ;
        RECT 111.510 23.445 111.680 33.485 ;
        RECT 113.090 23.445 113.260 33.485 ;
        RECT 114.670 23.445 114.840 33.485 ;
        RECT 116.250 23.445 116.420 33.485 ;
        RECT 117.830 23.445 118.000 33.485 ;
        RECT 119.410 23.445 119.580 33.485 ;
        RECT 124.920 32.020 125.250 33.000 ;
        RECT 123.380 31.845 124.210 31.935 ;
        RECT 124.520 31.845 124.850 31.850 ;
        RECT 123.380 31.615 124.850 31.845 ;
        RECT 123.380 31.415 124.210 31.615 ;
        RECT 124.520 31.610 124.850 31.615 ;
        RECT 125.020 31.805 125.250 32.020 ;
        RECT 126.580 32.765 126.910 32.990 ;
        RECT 126.580 32.205 127.290 32.765 ;
        RECT 126.580 32.010 126.910 32.205 ;
        RECT 126.180 31.805 126.510 31.840 ;
        RECT 125.020 31.615 126.510 31.805 ;
        RECT 125.020 31.420 125.250 31.615 ;
        RECT 126.180 31.600 126.510 31.615 ;
        RECT 124.920 30.790 125.250 31.420 ;
        RECT 126.680 31.410 126.910 32.010 ;
        RECT 126.580 30.780 126.910 31.410 ;
        RECT 125.750 29.875 127.830 30.195 ;
        RECT 125.750 29.795 126.820 29.875 ;
        RECT 127.310 29.795 127.830 29.875 ;
        RECT 125.750 29.620 125.990 29.795 ;
        RECT 125.745 29.270 125.995 29.620 ;
        RECT 126.175 29.100 126.815 29.170 ;
        RECT 125.405 28.930 126.815 29.100 ;
        RECT 125.405 28.750 125.575 28.930 ;
        RECT 126.175 28.840 126.815 28.930 ;
        RECT 124.620 28.420 125.575 28.750 ;
        RECT 125.745 28.410 125.995 28.760 ;
        RECT 125.750 28.235 125.990 28.410 ;
        RECT 125.740 27.775 125.990 28.235 ;
        RECT 124.635 27.545 126.845 27.775 ;
        RECT 124.635 27.445 125.615 27.545 ;
        RECT 126.215 27.445 126.845 27.545 ;
        RECT 23.390 23.060 23.890 23.230 ;
        RECT 24.180 23.060 24.680 23.230 ;
        RECT 24.970 23.060 25.470 23.230 ;
        RECT 25.760 23.060 26.260 23.230 ;
        RECT 26.550 23.060 27.050 23.230 ;
        RECT 27.340 23.060 27.840 23.230 ;
        RECT 28.130 23.060 28.630 23.230 ;
        RECT 28.920 23.060 29.420 23.230 ;
        RECT 29.710 23.060 30.210 23.230 ;
        RECT 30.500 23.060 31.000 23.230 ;
        RECT 31.290 23.060 31.790 23.230 ;
        RECT 32.080 23.060 32.580 23.230 ;
        RECT 32.870 23.060 33.370 23.230 ;
        RECT 33.660 23.060 34.160 23.230 ;
        RECT 34.450 23.060 34.950 23.230 ;
        RECT 35.240 23.060 35.740 23.230 ;
        RECT 36.030 23.060 36.530 23.230 ;
        RECT 36.820 23.060 37.320 23.230 ;
        RECT 105.420 23.060 105.920 23.230 ;
        RECT 106.210 23.060 106.710 23.230 ;
        RECT 107.000 23.060 107.500 23.230 ;
        RECT 107.790 23.060 108.290 23.230 ;
        RECT 108.580 23.060 109.080 23.230 ;
        RECT 109.370 23.060 109.870 23.230 ;
        RECT 110.160 23.060 110.660 23.230 ;
        RECT 110.950 23.060 111.450 23.230 ;
        RECT 111.740 23.060 112.240 23.230 ;
        RECT 112.530 23.060 113.030 23.230 ;
        RECT 113.320 23.060 113.820 23.230 ;
        RECT 114.110 23.060 114.610 23.230 ;
        RECT 114.900 23.060 115.400 23.230 ;
        RECT 115.690 23.060 116.190 23.230 ;
        RECT 116.480 23.060 116.980 23.230 ;
        RECT 117.270 23.060 117.770 23.230 ;
        RECT 118.060 23.060 118.560 23.230 ;
        RECT 118.850 23.060 119.350 23.230 ;
      LAYER met1 ;
        RECT 22.925 214.835 37.555 215.065 ;
        RECT 22.625 204.625 22.895 214.635 ;
        RECT 24.205 204.625 24.475 214.635 ;
        RECT 25.785 204.625 26.055 214.635 ;
        RECT 27.365 204.625 27.635 214.635 ;
        RECT 28.945 204.625 29.215 214.635 ;
        RECT 30.525 204.625 30.795 214.635 ;
        RECT 32.105 204.625 32.375 214.635 ;
        RECT 33.685 204.625 33.955 214.635 ;
        RECT 35.265 204.625 35.535 214.635 ;
        RECT 36.845 204.625 37.115 214.635 ;
        RECT 37.325 204.425 37.555 214.835 ;
        RECT 105.515 214.835 120.145 215.065 ;
        RECT 105.515 204.425 105.745 214.835 ;
        RECT 105.955 204.625 106.225 214.635 ;
        RECT 107.535 204.625 107.805 214.635 ;
        RECT 109.115 204.625 109.385 214.635 ;
        RECT 110.695 204.625 110.965 214.635 ;
        RECT 112.275 204.625 112.545 214.635 ;
        RECT 113.855 204.625 114.125 214.635 ;
        RECT 115.435 204.625 115.705 214.635 ;
        RECT 117.015 204.625 117.285 214.635 ;
        RECT 118.595 204.625 118.865 214.635 ;
        RECT 120.175 204.625 120.445 214.635 ;
        RECT 22.925 204.195 38.255 204.425 ;
        RECT 38.025 202.785 38.255 204.195 ;
        RECT 34.715 202.555 38.255 202.785 ;
        RECT 104.815 204.195 120.145 204.425 ;
        RECT 104.815 202.785 105.045 204.195 ;
        RECT 104.815 202.555 108.355 202.785 ;
        RECT 22.775 201.265 32.665 201.495 ;
        RECT 22.475 196.105 22.745 201.105 ;
        RECT 24.055 196.105 24.325 201.105 ;
        RECT 25.635 196.105 25.905 201.105 ;
        RECT 27.215 196.105 27.485 201.105 ;
        RECT 28.795 196.105 29.065 201.105 ;
        RECT 30.375 196.105 30.645 201.105 ;
        RECT 31.955 196.105 32.225 201.105 ;
        RECT 32.435 198.485 32.665 201.265 ;
        RECT 34.715 201.275 34.945 202.555 ;
        RECT 37.545 202.065 38.835 202.295 ;
        RECT 35.815 201.275 36.045 201.945 ;
        RECT 34.715 201.025 36.045 201.275 ;
        RECT 37.495 201.035 38.465 201.265 ;
        RECT 35.815 200.355 36.045 201.025 ;
        RECT 37.195 199.955 38.085 200.185 ;
        RECT 35.815 198.485 36.045 199.155 ;
        RECT 32.435 198.235 36.045 198.485 ;
        RECT 37.195 198.475 37.425 199.955 ;
        RECT 38.225 199.555 38.465 201.035 ;
        RECT 37.565 199.325 38.465 199.555 ;
        RECT 37.195 198.245 38.155 198.475 ;
        RECT 32.435 195.945 32.665 198.235 ;
        RECT 35.815 197.565 36.045 198.235 ;
        RECT 37.545 197.215 38.195 197.445 ;
        RECT 37.545 196.985 37.715 197.215 ;
        RECT 22.775 195.715 32.665 195.945 ;
        RECT 36.305 196.815 37.715 196.985 ;
        RECT 34.315 194.865 34.635 194.925 ;
        RECT 36.305 194.865 36.475 196.815 ;
        RECT 38.665 196.205 38.835 202.065 ;
        RECT 36.685 195.915 38.835 196.205 ;
        RECT 104.235 202.065 105.525 202.295 ;
        RECT 104.235 196.205 104.405 202.065 ;
        RECT 107.025 201.275 107.255 201.945 ;
        RECT 108.125 201.275 108.355 202.555 ;
        RECT 104.605 201.035 105.575 201.265 ;
        RECT 104.605 199.555 104.845 201.035 ;
        RECT 107.025 201.025 108.355 201.275 ;
        RECT 110.405 201.265 120.295 201.495 ;
        RECT 107.025 200.355 107.255 201.025 ;
        RECT 104.985 199.955 105.875 200.185 ;
        RECT 104.605 199.325 105.505 199.555 ;
        RECT 105.645 198.475 105.875 199.955 ;
        RECT 104.915 198.245 105.875 198.475 ;
        RECT 107.025 198.485 107.255 199.155 ;
        RECT 110.405 198.485 110.635 201.265 ;
        RECT 107.025 198.235 110.635 198.485 ;
        RECT 107.025 197.565 107.255 198.235 ;
        RECT 104.875 197.215 105.525 197.445 ;
        RECT 105.355 196.985 105.525 197.215 ;
        RECT 105.355 196.815 106.765 196.985 ;
        RECT 104.235 195.915 106.385 196.205 ;
        RECT 37.265 195.485 37.495 195.775 ;
        RECT 105.575 195.485 105.805 195.775 ;
        RECT 37.295 194.865 37.465 195.485 ;
        RECT 34.315 194.695 37.465 194.865 ;
        RECT 105.605 194.865 105.775 195.485 ;
        RECT 106.595 194.865 106.765 196.815 ;
        RECT 110.405 195.945 110.635 198.235 ;
        RECT 110.845 196.105 111.115 201.105 ;
        RECT 112.425 196.105 112.695 201.105 ;
        RECT 114.005 196.105 114.275 201.105 ;
        RECT 115.585 196.105 115.855 201.105 ;
        RECT 117.165 196.105 117.435 201.105 ;
        RECT 118.745 196.105 119.015 201.105 ;
        RECT 120.325 196.105 120.595 201.105 ;
        RECT 110.405 195.715 120.295 195.945 ;
        RECT 108.435 194.865 108.755 194.925 ;
        RECT 105.605 194.695 108.755 194.865 ;
        RECT 34.315 194.665 34.635 194.695 ;
        RECT 108.435 194.665 108.755 194.695 ;
        RECT 39.590 192.935 40.960 192.945 ;
        RECT 39.590 192.915 42.920 192.935 ;
        RECT 102.110 192.930 103.480 192.945 ;
        RECT 38.600 192.870 42.920 192.915 ;
        RECT 100.590 192.915 103.480 192.930 ;
        RECT 100.590 192.910 104.470 192.915 ;
        RECT 38.600 191.860 45.590 192.870 ;
        RECT 38.600 191.845 40.960 191.860 ;
        RECT 38.600 191.815 39.970 191.845 ;
        RECT 41.740 191.800 45.590 191.860 ;
        RECT 97.500 191.920 104.470 192.910 ;
        RECT 97.500 191.840 101.350 191.920 ;
        RECT 102.110 191.845 104.470 191.920 ;
        RECT 18.330 191.775 18.990 191.795 ;
        RECT 19.190 191.775 21.110 191.795 ;
        RECT 18.330 191.770 22.500 191.775 ;
        RECT 25.260 191.770 25.580 191.800 ;
        RECT 18.330 191.600 25.580 191.770 ;
        RECT 18.330 191.585 22.600 191.600 ;
        RECT 18.330 191.185 18.990 191.585 ;
        RECT 19.190 191.575 21.110 191.585 ;
        RECT 22.430 190.980 22.600 191.585 ;
        RECT 22.400 190.690 22.630 190.980 ;
        RECT 21.060 190.260 23.210 190.550 ;
        RECT 13.580 185.735 14.240 186.755 ;
        RECT 18.520 186.295 19.310 186.995 ;
        RECT 13.640 183.705 14.280 184.725 ;
        RECT 21.060 184.400 21.230 190.260 ;
        RECT 23.420 189.650 23.590 191.600 ;
        RECT 25.260 191.540 25.580 191.600 ;
        RECT 22.180 189.480 23.590 189.650 ;
        RECT 27.230 190.520 37.120 190.750 ;
        RECT 22.180 189.250 22.350 189.480 ;
        RECT 21.700 189.020 22.350 189.250 ;
        RECT 23.850 188.230 24.080 188.900 ;
        RECT 27.230 188.230 27.460 190.520 ;
        RECT 21.740 187.990 22.700 188.220 ;
        RECT 21.430 186.910 22.330 187.140 ;
        RECT 21.430 185.430 21.670 186.910 ;
        RECT 22.470 186.510 22.700 187.990 ;
        RECT 23.850 187.980 27.460 188.230 ;
        RECT 23.850 187.310 24.080 187.980 ;
        RECT 21.810 186.280 22.700 186.510 ;
        RECT 23.850 185.440 24.080 186.110 ;
        RECT 21.430 185.200 22.400 185.430 ;
        RECT 23.850 185.190 25.180 185.440 ;
        RECT 23.850 184.520 24.080 185.190 ;
        RECT 21.060 184.170 22.350 184.400 ;
        RECT 24.950 183.910 25.180 185.190 ;
        RECT 27.230 185.200 27.460 187.980 ;
        RECT 27.670 185.360 27.940 190.360 ;
        RECT 29.250 185.360 29.520 190.360 ;
        RECT 30.830 185.360 31.100 190.360 ;
        RECT 32.410 185.360 32.680 190.360 ;
        RECT 33.990 185.360 34.260 190.360 ;
        RECT 35.570 185.360 35.840 190.360 ;
        RECT 37.150 185.360 37.420 190.360 ;
        RECT 27.230 184.970 37.120 185.200 ;
        RECT 42.840 183.970 44.880 191.800 ;
        RECT 98.210 184.010 100.250 191.840 ;
        RECT 103.100 191.815 104.470 191.845 ;
        RECT 117.490 191.770 117.810 191.800 ;
        RECT 121.960 191.775 123.880 191.795 ;
        RECT 124.080 191.775 124.740 191.795 ;
        RECT 120.570 191.770 124.740 191.775 ;
        RECT 117.490 191.600 124.740 191.770 ;
        RECT 117.490 191.540 117.810 191.600 ;
        RECT 105.950 190.520 115.840 190.750 ;
        RECT 105.650 185.360 105.920 190.360 ;
        RECT 107.230 185.360 107.500 190.360 ;
        RECT 108.810 185.360 109.080 190.360 ;
        RECT 110.390 185.360 110.660 190.360 ;
        RECT 111.970 185.360 112.240 190.360 ;
        RECT 113.550 185.360 113.820 190.360 ;
        RECT 115.130 185.360 115.400 190.360 ;
        RECT 115.610 188.230 115.840 190.520 ;
        RECT 119.480 189.650 119.650 191.600 ;
        RECT 120.470 191.585 124.740 191.600 ;
        RECT 120.470 190.980 120.640 191.585 ;
        RECT 121.960 191.575 123.880 191.585 ;
        RECT 124.080 191.185 124.740 191.585 ;
        RECT 120.440 190.690 120.670 190.980 ;
        RECT 119.860 190.260 122.010 190.550 ;
        RECT 119.480 189.480 120.890 189.650 ;
        RECT 120.720 189.250 120.890 189.480 ;
        RECT 120.720 189.020 121.370 189.250 ;
        RECT 118.990 188.230 119.220 188.900 ;
        RECT 115.610 187.980 119.220 188.230 ;
        RECT 115.610 185.200 115.840 187.980 ;
        RECT 118.990 187.310 119.220 187.980 ;
        RECT 120.370 187.990 121.330 188.220 ;
        RECT 120.370 186.510 120.600 187.990 ;
        RECT 120.740 186.910 121.640 187.140 ;
        RECT 120.370 186.280 121.260 186.510 ;
        RECT 118.990 185.440 119.220 186.110 ;
        RECT 105.950 184.970 115.840 185.200 ;
        RECT 117.890 185.190 119.220 185.440 ;
        RECT 121.400 185.430 121.640 186.910 ;
        RECT 120.670 185.200 121.640 185.430 ;
        RECT 21.640 183.680 25.180 183.910 ;
        RECT 117.890 183.910 118.120 185.190 ;
        RECT 118.990 184.520 119.220 185.190 ;
        RECT 121.840 184.400 122.010 190.260 ;
        RECT 123.760 186.295 124.550 186.995 ;
        RECT 128.830 185.735 129.490 186.755 ;
        RECT 120.720 184.170 122.010 184.400 ;
        RECT 117.890 183.680 121.430 183.910 ;
        RECT 128.790 183.705 129.430 184.725 ;
        RECT 21.640 182.270 21.870 183.680 ;
        RECT 121.200 182.270 121.430 183.680 ;
        RECT 21.640 182.040 36.970 182.270 ;
        RECT 106.100 182.040 121.430 182.270 ;
        RECT 15.060 181.125 15.790 181.155 ;
        RECT 15.060 181.055 15.850 181.125 ;
        RECT 15.040 180.635 15.850 181.055 ;
        RECT 15.060 180.585 15.850 180.635 ;
        RECT 15.060 180.555 15.790 180.585 ;
        RECT 18.160 179.755 19.100 180.345 ;
        RECT 16.840 178.495 17.660 178.525 ;
        RECT 14.610 178.415 14.960 178.465 ;
        RECT 14.350 178.385 14.960 178.415 ;
        RECT 14.320 178.215 14.980 178.385 ;
        RECT 14.320 177.785 14.960 178.215 ;
        RECT 16.840 178.025 17.680 178.495 ;
        RECT 16.840 177.995 17.660 178.025 ;
        RECT 14.340 177.745 14.960 177.785 ;
        RECT 17.130 177.515 17.470 177.995 ;
        RECT 17.120 177.355 17.470 177.515 ;
        RECT 17.110 177.275 17.470 177.355 ;
        RECT 17.110 177.085 17.460 177.275 ;
        RECT 17.110 176.965 17.510 177.085 ;
        RECT 17.140 176.845 17.510 176.965 ;
        RECT 17.140 176.785 17.490 176.845 ;
        RECT 22.340 171.630 22.570 182.040 ;
        RECT 22.780 171.830 23.050 181.840 ;
        RECT 24.360 171.830 24.630 181.840 ;
        RECT 25.940 171.830 26.210 181.840 ;
        RECT 27.520 171.830 27.790 181.840 ;
        RECT 29.100 171.830 29.370 181.840 ;
        RECT 30.680 171.830 30.950 181.840 ;
        RECT 32.260 171.830 32.530 181.840 ;
        RECT 33.840 171.830 34.110 181.840 ;
        RECT 35.420 171.830 35.690 181.840 ;
        RECT 37.000 171.830 37.270 181.840 ;
        RECT 105.800 171.830 106.070 181.840 ;
        RECT 107.380 171.830 107.650 181.840 ;
        RECT 108.960 171.830 109.230 181.840 ;
        RECT 110.540 171.830 110.810 181.840 ;
        RECT 112.120 171.830 112.390 181.840 ;
        RECT 113.700 171.830 113.970 181.840 ;
        RECT 115.280 171.830 115.550 181.840 ;
        RECT 116.860 171.830 117.130 181.840 ;
        RECT 118.440 171.830 118.710 181.840 ;
        RECT 120.020 171.830 120.290 181.840 ;
        RECT 120.500 171.630 120.730 182.040 ;
        RECT 127.280 181.125 128.010 181.155 ;
        RECT 127.220 181.055 128.010 181.125 ;
        RECT 127.220 180.635 128.030 181.055 ;
        RECT 127.220 180.585 128.010 180.635 ;
        RECT 127.280 180.555 128.010 180.585 ;
        RECT 123.970 179.755 124.910 180.345 ;
        RECT 125.410 178.495 126.230 178.525 ;
        RECT 125.390 178.025 126.230 178.495 ;
        RECT 128.110 178.415 128.460 178.465 ;
        RECT 128.110 178.385 128.720 178.415 ;
        RECT 128.090 178.215 128.750 178.385 ;
        RECT 125.410 177.995 126.230 178.025 ;
        RECT 125.600 177.515 125.940 177.995 ;
        RECT 128.110 177.785 128.750 178.215 ;
        RECT 128.110 177.745 128.730 177.785 ;
        RECT 125.600 177.355 125.950 177.515 ;
        RECT 125.600 177.275 125.960 177.355 ;
        RECT 125.610 177.085 125.960 177.275 ;
        RECT 125.560 176.965 125.960 177.085 ;
        RECT 125.560 176.845 125.930 176.965 ;
        RECT 125.580 176.785 125.930 176.845 ;
        RECT 22.340 171.400 36.970 171.630 ;
        RECT 106.100 171.400 120.730 171.630 ;
        RECT 22.925 165.265 37.555 165.495 ;
        RECT 22.625 155.055 22.895 165.065 ;
        RECT 24.205 155.055 24.475 165.065 ;
        RECT 25.785 155.055 26.055 165.065 ;
        RECT 27.365 155.055 27.635 165.065 ;
        RECT 28.945 155.055 29.215 165.065 ;
        RECT 30.525 155.055 30.795 165.065 ;
        RECT 32.105 155.055 32.375 165.065 ;
        RECT 33.685 155.055 33.955 165.065 ;
        RECT 35.265 155.055 35.535 165.065 ;
        RECT 36.845 155.055 37.115 165.065 ;
        RECT 37.325 154.855 37.555 165.265 ;
        RECT 105.515 165.265 120.145 165.495 ;
        RECT 105.515 154.855 105.745 165.265 ;
        RECT 105.955 155.055 106.225 165.065 ;
        RECT 107.535 155.055 107.805 165.065 ;
        RECT 109.115 155.055 109.385 165.065 ;
        RECT 110.695 155.055 110.965 165.065 ;
        RECT 112.275 155.055 112.545 165.065 ;
        RECT 113.855 155.055 114.125 165.065 ;
        RECT 115.435 155.055 115.705 165.065 ;
        RECT 117.015 155.055 117.285 165.065 ;
        RECT 118.595 155.055 118.865 165.065 ;
        RECT 120.175 155.055 120.445 165.065 ;
        RECT 22.925 154.625 38.255 154.855 ;
        RECT 38.025 153.215 38.255 154.625 ;
        RECT 34.715 152.985 38.255 153.215 ;
        RECT 104.815 154.625 120.145 154.855 ;
        RECT 104.815 153.215 105.045 154.625 ;
        RECT 104.815 152.985 108.355 153.215 ;
        RECT 22.775 151.695 32.665 151.925 ;
        RECT 22.475 146.535 22.745 151.535 ;
        RECT 24.055 146.535 24.325 151.535 ;
        RECT 25.635 146.535 25.905 151.535 ;
        RECT 27.215 146.535 27.485 151.535 ;
        RECT 28.795 146.535 29.065 151.535 ;
        RECT 30.375 146.535 30.645 151.535 ;
        RECT 31.955 146.535 32.225 151.535 ;
        RECT 32.435 148.915 32.665 151.695 ;
        RECT 34.715 151.705 34.945 152.985 ;
        RECT 37.545 152.495 38.835 152.725 ;
        RECT 35.815 151.705 36.045 152.375 ;
        RECT 34.715 151.455 36.045 151.705 ;
        RECT 37.495 151.465 38.465 151.695 ;
        RECT 35.815 150.785 36.045 151.455 ;
        RECT 37.195 150.385 38.085 150.615 ;
        RECT 35.815 148.915 36.045 149.585 ;
        RECT 32.435 148.665 36.045 148.915 ;
        RECT 37.195 148.905 37.425 150.385 ;
        RECT 38.225 149.985 38.465 151.465 ;
        RECT 37.565 149.755 38.465 149.985 ;
        RECT 37.195 148.675 38.155 148.905 ;
        RECT 32.435 146.375 32.665 148.665 ;
        RECT 35.815 147.995 36.045 148.665 ;
        RECT 37.545 147.645 38.195 147.875 ;
        RECT 37.545 147.415 37.715 147.645 ;
        RECT 22.775 146.145 32.665 146.375 ;
        RECT 36.305 147.245 37.715 147.415 ;
        RECT 34.315 145.295 34.635 145.355 ;
        RECT 36.305 145.295 36.475 147.245 ;
        RECT 38.665 146.635 38.835 152.495 ;
        RECT 36.685 146.345 38.835 146.635 ;
        RECT 104.235 152.495 105.525 152.725 ;
        RECT 104.235 146.635 104.405 152.495 ;
        RECT 107.025 151.705 107.255 152.375 ;
        RECT 108.125 151.705 108.355 152.985 ;
        RECT 104.605 151.465 105.575 151.695 ;
        RECT 104.605 149.985 104.845 151.465 ;
        RECT 107.025 151.455 108.355 151.705 ;
        RECT 110.405 151.695 120.295 151.925 ;
        RECT 107.025 150.785 107.255 151.455 ;
        RECT 104.985 150.385 105.875 150.615 ;
        RECT 104.605 149.755 105.505 149.985 ;
        RECT 105.645 148.905 105.875 150.385 ;
        RECT 104.915 148.675 105.875 148.905 ;
        RECT 107.025 148.915 107.255 149.585 ;
        RECT 110.405 148.915 110.635 151.695 ;
        RECT 107.025 148.665 110.635 148.915 ;
        RECT 107.025 147.995 107.255 148.665 ;
        RECT 104.875 147.645 105.525 147.875 ;
        RECT 105.355 147.415 105.525 147.645 ;
        RECT 105.355 147.245 106.765 147.415 ;
        RECT 104.235 146.345 106.385 146.635 ;
        RECT 37.265 145.915 37.495 146.205 ;
        RECT 105.575 145.915 105.805 146.205 ;
        RECT 37.295 145.295 37.465 145.915 ;
        RECT 34.315 145.125 37.465 145.295 ;
        RECT 105.605 145.295 105.775 145.915 ;
        RECT 106.595 145.295 106.765 147.245 ;
        RECT 110.405 146.375 110.635 148.665 ;
        RECT 110.845 146.535 111.115 151.535 ;
        RECT 112.425 146.535 112.695 151.535 ;
        RECT 114.005 146.535 114.275 151.535 ;
        RECT 115.585 146.535 115.855 151.535 ;
        RECT 117.165 146.535 117.435 151.535 ;
        RECT 118.745 146.535 119.015 151.535 ;
        RECT 120.325 146.535 120.595 151.535 ;
        RECT 110.405 146.145 120.295 146.375 ;
        RECT 108.435 145.295 108.755 145.355 ;
        RECT 105.605 145.125 108.755 145.295 ;
        RECT 34.315 145.095 34.635 145.125 ;
        RECT 108.435 145.095 108.755 145.125 ;
        RECT 39.590 143.345 42.540 143.375 ;
        RECT 102.110 143.355 103.480 143.375 ;
        RECT 101.940 143.350 103.480 143.355 ;
        RECT 38.600 143.340 42.540 143.345 ;
        RECT 100.170 143.345 103.480 143.350 ;
        RECT 38.600 142.300 45.640 143.340 ;
        RECT 100.170 143.300 104.470 143.345 ;
        RECT 38.600 142.275 40.960 142.300 ;
        RECT 38.600 142.245 39.970 142.275 ;
        RECT 41.790 142.270 45.640 142.300 ;
        RECT 97.370 142.340 104.470 143.300 ;
        RECT 18.330 142.205 18.990 142.225 ;
        RECT 19.190 142.205 21.110 142.225 ;
        RECT 18.330 142.200 22.500 142.205 ;
        RECT 25.260 142.200 25.580 142.230 ;
        RECT 18.330 142.030 25.580 142.200 ;
        RECT 18.330 142.015 22.600 142.030 ;
        RECT 18.330 141.615 18.990 142.015 ;
        RECT 19.190 142.005 21.110 142.015 ;
        RECT 22.430 141.410 22.600 142.015 ;
        RECT 22.400 141.120 22.630 141.410 ;
        RECT 21.060 140.690 23.210 140.980 ;
        RECT 13.580 136.165 14.240 137.185 ;
        RECT 18.520 136.725 19.310 137.425 ;
        RECT 13.640 134.135 14.280 135.155 ;
        RECT 21.060 134.830 21.230 140.690 ;
        RECT 23.420 140.080 23.590 142.030 ;
        RECT 25.260 141.970 25.580 142.030 ;
        RECT 22.180 139.910 23.590 140.080 ;
        RECT 27.230 140.950 37.120 141.180 ;
        RECT 22.180 139.680 22.350 139.910 ;
        RECT 21.700 139.450 22.350 139.680 ;
        RECT 23.850 138.660 24.080 139.330 ;
        RECT 27.230 138.660 27.460 140.950 ;
        RECT 21.740 138.420 22.700 138.650 ;
        RECT 21.430 137.340 22.330 137.570 ;
        RECT 21.430 135.860 21.670 137.340 ;
        RECT 22.470 136.940 22.700 138.420 ;
        RECT 23.850 138.410 27.460 138.660 ;
        RECT 23.850 137.740 24.080 138.410 ;
        RECT 21.810 136.710 22.700 136.940 ;
        RECT 23.850 135.870 24.080 136.540 ;
        RECT 21.430 135.630 22.400 135.860 ;
        RECT 23.850 135.620 25.180 135.870 ;
        RECT 23.850 134.950 24.080 135.620 ;
        RECT 21.060 134.600 22.350 134.830 ;
        RECT 24.950 134.340 25.180 135.620 ;
        RECT 27.230 135.630 27.460 138.410 ;
        RECT 27.670 135.790 27.940 140.790 ;
        RECT 29.250 135.790 29.520 140.790 ;
        RECT 30.830 135.790 31.100 140.790 ;
        RECT 32.410 135.790 32.680 140.790 ;
        RECT 33.990 135.790 34.260 140.790 ;
        RECT 35.570 135.790 35.840 140.790 ;
        RECT 37.150 135.790 37.420 140.790 ;
        RECT 27.230 135.400 37.120 135.630 ;
        RECT 42.890 134.440 44.930 142.270 ;
        RECT 97.370 142.230 101.220 142.340 ;
        RECT 102.110 142.275 104.470 142.340 ;
        RECT 103.100 142.245 104.470 142.275 ;
        RECT 98.080 134.400 100.120 142.230 ;
        RECT 117.490 142.200 117.810 142.230 ;
        RECT 121.960 142.205 123.880 142.225 ;
        RECT 124.080 142.205 124.740 142.225 ;
        RECT 120.570 142.200 124.740 142.205 ;
        RECT 117.490 142.030 124.740 142.200 ;
        RECT 117.490 141.970 117.810 142.030 ;
        RECT 105.950 140.950 115.840 141.180 ;
        RECT 105.650 135.790 105.920 140.790 ;
        RECT 107.230 135.790 107.500 140.790 ;
        RECT 108.810 135.790 109.080 140.790 ;
        RECT 110.390 135.790 110.660 140.790 ;
        RECT 111.970 135.790 112.240 140.790 ;
        RECT 113.550 135.790 113.820 140.790 ;
        RECT 115.130 135.790 115.400 140.790 ;
        RECT 115.610 138.660 115.840 140.950 ;
        RECT 119.480 140.080 119.650 142.030 ;
        RECT 120.470 142.015 124.740 142.030 ;
        RECT 120.470 141.410 120.640 142.015 ;
        RECT 121.960 142.005 123.880 142.015 ;
        RECT 124.080 141.615 124.740 142.015 ;
        RECT 120.440 141.120 120.670 141.410 ;
        RECT 119.860 140.690 122.010 140.980 ;
        RECT 119.480 139.910 120.890 140.080 ;
        RECT 120.720 139.680 120.890 139.910 ;
        RECT 120.720 139.450 121.370 139.680 ;
        RECT 118.990 138.660 119.220 139.330 ;
        RECT 115.610 138.410 119.220 138.660 ;
        RECT 115.610 135.630 115.840 138.410 ;
        RECT 118.990 137.740 119.220 138.410 ;
        RECT 120.370 138.420 121.330 138.650 ;
        RECT 120.370 136.940 120.600 138.420 ;
        RECT 120.740 137.340 121.640 137.570 ;
        RECT 120.370 136.710 121.260 136.940 ;
        RECT 118.990 135.870 119.220 136.540 ;
        RECT 105.950 135.400 115.840 135.630 ;
        RECT 117.890 135.620 119.220 135.870 ;
        RECT 121.400 135.860 121.640 137.340 ;
        RECT 120.670 135.630 121.640 135.860 ;
        RECT 21.640 134.110 25.180 134.340 ;
        RECT 117.890 134.340 118.120 135.620 ;
        RECT 118.990 134.950 119.220 135.620 ;
        RECT 121.840 134.830 122.010 140.690 ;
        RECT 123.760 136.725 124.550 137.425 ;
        RECT 128.830 136.165 129.490 137.185 ;
        RECT 120.720 134.600 122.010 134.830 ;
        RECT 117.890 134.110 121.430 134.340 ;
        RECT 128.790 134.135 129.430 135.155 ;
        RECT 21.640 132.700 21.870 134.110 ;
        RECT 121.200 132.700 121.430 134.110 ;
        RECT 21.640 132.470 36.970 132.700 ;
        RECT 106.100 132.470 121.430 132.700 ;
        RECT 15.060 131.555 15.790 131.585 ;
        RECT 15.060 131.485 15.850 131.555 ;
        RECT 15.040 131.065 15.850 131.485 ;
        RECT 15.060 131.015 15.850 131.065 ;
        RECT 15.060 130.985 15.790 131.015 ;
        RECT 18.160 130.185 19.100 130.775 ;
        RECT 16.840 128.925 17.660 128.955 ;
        RECT 14.610 128.845 14.960 128.895 ;
        RECT 14.350 128.815 14.960 128.845 ;
        RECT 14.320 128.645 14.980 128.815 ;
        RECT 14.320 128.215 14.960 128.645 ;
        RECT 16.840 128.455 17.680 128.925 ;
        RECT 16.840 128.425 17.660 128.455 ;
        RECT 14.340 128.175 14.960 128.215 ;
        RECT 17.130 127.945 17.470 128.425 ;
        RECT 17.120 127.785 17.470 127.945 ;
        RECT 17.110 127.705 17.470 127.785 ;
        RECT 17.110 127.515 17.460 127.705 ;
        RECT 17.110 127.395 17.510 127.515 ;
        RECT 17.140 127.275 17.510 127.395 ;
        RECT 17.140 127.215 17.490 127.275 ;
        RECT 22.340 122.060 22.570 132.470 ;
        RECT 22.780 122.260 23.050 132.270 ;
        RECT 24.360 122.260 24.630 132.270 ;
        RECT 25.940 122.260 26.210 132.270 ;
        RECT 27.520 122.260 27.790 132.270 ;
        RECT 29.100 122.260 29.370 132.270 ;
        RECT 30.680 122.260 30.950 132.270 ;
        RECT 32.260 122.260 32.530 132.270 ;
        RECT 33.840 122.260 34.110 132.270 ;
        RECT 35.420 122.260 35.690 132.270 ;
        RECT 37.000 122.260 37.270 132.270 ;
        RECT 105.800 122.260 106.070 132.270 ;
        RECT 107.380 122.260 107.650 132.270 ;
        RECT 108.960 122.260 109.230 132.270 ;
        RECT 110.540 122.260 110.810 132.270 ;
        RECT 112.120 122.260 112.390 132.270 ;
        RECT 113.700 122.260 113.970 132.270 ;
        RECT 115.280 122.260 115.550 132.270 ;
        RECT 116.860 122.260 117.130 132.270 ;
        RECT 118.440 122.260 118.710 132.270 ;
        RECT 120.020 122.260 120.290 132.270 ;
        RECT 120.500 122.060 120.730 132.470 ;
        RECT 127.280 131.555 128.010 131.585 ;
        RECT 127.220 131.485 128.010 131.555 ;
        RECT 127.220 131.065 128.030 131.485 ;
        RECT 127.220 131.015 128.010 131.065 ;
        RECT 127.280 130.985 128.010 131.015 ;
        RECT 123.970 130.185 124.910 130.775 ;
        RECT 125.410 128.925 126.230 128.955 ;
        RECT 125.390 128.455 126.230 128.925 ;
        RECT 128.110 128.845 128.460 128.895 ;
        RECT 128.110 128.815 128.720 128.845 ;
        RECT 128.090 128.645 128.750 128.815 ;
        RECT 125.410 128.425 126.230 128.455 ;
        RECT 125.600 127.945 125.940 128.425 ;
        RECT 128.110 128.215 128.750 128.645 ;
        RECT 128.110 128.175 128.730 128.215 ;
        RECT 125.600 127.785 125.950 127.945 ;
        RECT 125.600 127.705 125.960 127.785 ;
        RECT 125.610 127.515 125.960 127.705 ;
        RECT 125.560 127.395 125.960 127.515 ;
        RECT 125.560 127.275 125.930 127.395 ;
        RECT 125.580 127.215 125.930 127.275 ;
        RECT 22.340 121.830 36.970 122.060 ;
        RECT 106.100 121.830 120.730 122.060 ;
        RECT 23.585 117.035 38.215 117.265 ;
        RECT 23.285 106.825 23.555 116.835 ;
        RECT 24.865 106.825 25.135 116.835 ;
        RECT 26.445 106.825 26.715 116.835 ;
        RECT 28.025 106.825 28.295 116.835 ;
        RECT 29.605 106.825 29.875 116.835 ;
        RECT 31.185 106.825 31.455 116.835 ;
        RECT 32.765 106.825 33.035 116.835 ;
        RECT 34.345 106.825 34.615 116.835 ;
        RECT 35.925 106.825 36.195 116.835 ;
        RECT 37.505 106.825 37.775 116.835 ;
        RECT 37.985 106.625 38.215 117.035 ;
        RECT 105.515 116.365 120.145 116.595 ;
        RECT 23.585 106.395 38.915 106.625 ;
        RECT 38.685 104.985 38.915 106.395 ;
        RECT 105.515 105.955 105.745 116.365 ;
        RECT 105.955 106.155 106.225 116.165 ;
        RECT 107.535 106.155 107.805 116.165 ;
        RECT 109.115 106.155 109.385 116.165 ;
        RECT 110.695 106.155 110.965 116.165 ;
        RECT 112.275 106.155 112.545 116.165 ;
        RECT 113.855 106.155 114.125 116.165 ;
        RECT 115.435 106.155 115.705 116.165 ;
        RECT 117.015 106.155 117.285 116.165 ;
        RECT 118.595 106.155 118.865 116.165 ;
        RECT 120.175 106.155 120.445 116.165 ;
        RECT 35.375 104.755 38.915 104.985 ;
        RECT 104.815 105.725 120.145 105.955 ;
        RECT 23.435 103.465 33.325 103.695 ;
        RECT 23.135 98.305 23.405 103.305 ;
        RECT 24.715 98.305 24.985 103.305 ;
        RECT 26.295 98.305 26.565 103.305 ;
        RECT 27.875 98.305 28.145 103.305 ;
        RECT 29.455 98.305 29.725 103.305 ;
        RECT 31.035 98.305 31.305 103.305 ;
        RECT 32.615 98.305 32.885 103.305 ;
        RECT 33.095 100.685 33.325 103.465 ;
        RECT 35.375 103.475 35.605 104.755 ;
        RECT 38.205 104.265 39.495 104.495 ;
        RECT 36.475 103.475 36.705 104.145 ;
        RECT 35.375 103.225 36.705 103.475 ;
        RECT 38.155 103.235 39.125 103.465 ;
        RECT 36.475 102.555 36.705 103.225 ;
        RECT 37.855 102.155 38.745 102.385 ;
        RECT 36.475 100.685 36.705 101.355 ;
        RECT 33.095 100.435 36.705 100.685 ;
        RECT 37.855 100.675 38.085 102.155 ;
        RECT 38.885 101.755 39.125 103.235 ;
        RECT 38.225 101.525 39.125 101.755 ;
        RECT 37.855 100.445 38.815 100.675 ;
        RECT 33.095 98.145 33.325 100.435 ;
        RECT 36.475 99.765 36.705 100.435 ;
        RECT 38.205 99.415 38.855 99.645 ;
        RECT 38.205 99.185 38.375 99.415 ;
        RECT 23.435 97.915 33.325 98.145 ;
        RECT 36.965 99.015 38.375 99.185 ;
        RECT 34.975 97.065 35.295 97.125 ;
        RECT 36.965 97.065 37.135 99.015 ;
        RECT 39.325 98.405 39.495 104.265 ;
        RECT 104.815 104.315 105.045 105.725 ;
        RECT 104.815 104.085 108.355 104.315 ;
        RECT 37.345 98.115 39.495 98.405 ;
        RECT 104.235 103.595 105.525 103.825 ;
        RECT 37.925 97.685 38.155 97.975 ;
        RECT 104.235 97.735 104.405 103.595 ;
        RECT 107.025 102.805 107.255 103.475 ;
        RECT 108.125 102.805 108.355 104.085 ;
        RECT 104.605 102.565 105.575 102.795 ;
        RECT 104.605 101.085 104.845 102.565 ;
        RECT 107.025 102.555 108.355 102.805 ;
        RECT 110.405 102.795 120.295 103.025 ;
        RECT 107.025 101.885 107.255 102.555 ;
        RECT 104.985 101.485 105.875 101.715 ;
        RECT 104.605 100.855 105.505 101.085 ;
        RECT 105.645 100.005 105.875 101.485 ;
        RECT 104.915 99.775 105.875 100.005 ;
        RECT 107.025 100.015 107.255 100.685 ;
        RECT 110.405 100.015 110.635 102.795 ;
        RECT 107.025 99.765 110.635 100.015 ;
        RECT 107.025 99.095 107.255 99.765 ;
        RECT 104.875 98.745 105.525 98.975 ;
        RECT 105.355 98.515 105.525 98.745 ;
        RECT 105.355 98.345 106.765 98.515 ;
        RECT 37.955 97.065 38.125 97.685 ;
        RECT 104.235 97.445 106.385 97.735 ;
        RECT 34.975 96.895 38.125 97.065 ;
        RECT 105.575 97.015 105.805 97.305 ;
        RECT 34.975 96.865 35.295 96.895 ;
        RECT 105.605 96.395 105.775 97.015 ;
        RECT 106.595 96.395 106.765 98.345 ;
        RECT 110.405 97.475 110.635 99.765 ;
        RECT 110.845 97.635 111.115 102.635 ;
        RECT 112.425 97.635 112.695 102.635 ;
        RECT 114.005 97.635 114.275 102.635 ;
        RECT 115.585 97.635 115.855 102.635 ;
        RECT 117.165 97.635 117.435 102.635 ;
        RECT 118.745 97.635 119.015 102.635 ;
        RECT 120.325 97.635 120.595 102.635 ;
        RECT 110.405 97.245 120.295 97.475 ;
        RECT 108.435 96.395 108.755 96.455 ;
        RECT 105.605 96.225 108.755 96.395 ;
        RECT 108.435 96.195 108.755 96.225 ;
        RECT 41.570 95.150 42.610 95.180 ;
        RECT 41.570 95.145 46.140 95.150 ;
        RECT 40.250 95.115 46.140 95.145 ;
        RECT 39.260 94.080 46.140 95.115 ;
        RECT 102.110 94.455 103.480 94.475 ;
        RECT 101.940 94.445 103.480 94.455 ;
        RECT 101.940 94.390 104.470 94.445 ;
        RECT 99.970 94.360 104.470 94.390 ;
        RECT 39.260 94.070 42.610 94.080 ;
        RECT 39.260 94.045 41.620 94.070 ;
        RECT 39.260 94.015 40.630 94.045 ;
        RECT 18.990 93.975 19.650 93.995 ;
        RECT 19.850 93.975 21.770 93.995 ;
        RECT 18.990 93.970 23.160 93.975 ;
        RECT 25.920 93.970 26.240 94.000 ;
        RECT 18.990 93.800 26.240 93.970 ;
        RECT 18.990 93.785 23.260 93.800 ;
        RECT 18.990 93.385 19.650 93.785 ;
        RECT 19.850 93.775 21.770 93.785 ;
        RECT 23.090 93.180 23.260 93.785 ;
        RECT 23.060 92.890 23.290 93.180 ;
        RECT 21.720 92.460 23.870 92.750 ;
        RECT 14.240 87.935 14.900 88.955 ;
        RECT 19.180 88.495 19.970 89.195 ;
        RECT 14.300 85.905 14.940 86.925 ;
        RECT 21.720 86.600 21.890 92.460 ;
        RECT 24.080 91.850 24.250 93.800 ;
        RECT 25.920 93.740 26.240 93.800 ;
        RECT 22.840 91.680 24.250 91.850 ;
        RECT 27.890 92.720 37.780 92.950 ;
        RECT 22.840 91.450 23.010 91.680 ;
        RECT 22.360 91.220 23.010 91.450 ;
        RECT 24.510 90.430 24.740 91.100 ;
        RECT 27.890 90.430 28.120 92.720 ;
        RECT 22.400 90.190 23.360 90.420 ;
        RECT 22.090 89.110 22.990 89.340 ;
        RECT 22.090 87.630 22.330 89.110 ;
        RECT 23.130 88.710 23.360 90.190 ;
        RECT 24.510 90.180 28.120 90.430 ;
        RECT 24.510 89.510 24.740 90.180 ;
        RECT 22.470 88.480 23.360 88.710 ;
        RECT 24.510 87.640 24.740 88.310 ;
        RECT 22.090 87.400 23.060 87.630 ;
        RECT 24.510 87.390 25.840 87.640 ;
        RECT 24.510 86.720 24.740 87.390 ;
        RECT 21.720 86.370 23.010 86.600 ;
        RECT 25.610 86.110 25.840 87.390 ;
        RECT 27.890 87.400 28.120 90.180 ;
        RECT 28.330 87.560 28.600 92.560 ;
        RECT 29.910 87.560 30.180 92.560 ;
        RECT 31.490 87.560 31.760 92.560 ;
        RECT 33.070 87.560 33.340 92.560 ;
        RECT 34.650 87.560 34.920 92.560 ;
        RECT 36.230 87.560 36.500 92.560 ;
        RECT 37.810 87.560 38.080 92.560 ;
        RECT 27.890 87.170 37.780 87.400 ;
        RECT 43.390 86.250 45.430 94.080 ;
        RECT 97.460 93.380 104.470 94.360 ;
        RECT 97.460 93.290 101.310 93.380 ;
        RECT 102.110 93.375 104.470 93.380 ;
        RECT 103.100 93.345 104.470 93.375 ;
        RECT 117.490 93.300 117.810 93.330 ;
        RECT 121.960 93.305 123.880 93.325 ;
        RECT 124.080 93.305 124.740 93.325 ;
        RECT 120.570 93.300 124.740 93.305 ;
        RECT 22.300 85.880 25.840 86.110 ;
        RECT 22.300 84.470 22.530 85.880 ;
        RECT 98.170 85.460 100.210 93.290 ;
        RECT 117.490 93.130 124.740 93.300 ;
        RECT 117.490 93.070 117.810 93.130 ;
        RECT 105.950 92.050 115.840 92.280 ;
        RECT 105.650 86.890 105.920 91.890 ;
        RECT 107.230 86.890 107.500 91.890 ;
        RECT 108.810 86.890 109.080 91.890 ;
        RECT 110.390 86.890 110.660 91.890 ;
        RECT 111.970 86.890 112.240 91.890 ;
        RECT 113.550 86.890 113.820 91.890 ;
        RECT 115.130 86.890 115.400 91.890 ;
        RECT 115.610 89.760 115.840 92.050 ;
        RECT 119.480 91.180 119.650 93.130 ;
        RECT 120.470 93.115 124.740 93.130 ;
        RECT 120.470 92.510 120.640 93.115 ;
        RECT 121.960 93.105 123.880 93.115 ;
        RECT 124.080 92.715 124.740 93.115 ;
        RECT 120.440 92.220 120.670 92.510 ;
        RECT 119.860 91.790 122.010 92.080 ;
        RECT 119.480 91.010 120.890 91.180 ;
        RECT 120.720 90.780 120.890 91.010 ;
        RECT 120.720 90.550 121.370 90.780 ;
        RECT 118.990 89.760 119.220 90.430 ;
        RECT 115.610 89.510 119.220 89.760 ;
        RECT 115.610 86.730 115.840 89.510 ;
        RECT 118.990 88.840 119.220 89.510 ;
        RECT 120.370 89.520 121.330 89.750 ;
        RECT 120.370 88.040 120.600 89.520 ;
        RECT 120.740 88.440 121.640 88.670 ;
        RECT 120.370 87.810 121.260 88.040 ;
        RECT 118.990 86.970 119.220 87.640 ;
        RECT 105.950 86.500 115.840 86.730 ;
        RECT 117.890 86.720 119.220 86.970 ;
        RECT 121.400 86.960 121.640 88.440 ;
        RECT 120.670 86.730 121.640 86.960 ;
        RECT 117.890 85.440 118.120 86.720 ;
        RECT 118.990 86.050 119.220 86.720 ;
        RECT 121.840 85.930 122.010 91.790 ;
        RECT 123.760 87.825 124.550 88.525 ;
        RECT 128.830 87.265 129.490 88.285 ;
        RECT 120.720 85.700 122.010 85.930 ;
        RECT 117.890 85.210 121.430 85.440 ;
        RECT 128.790 85.235 129.430 86.255 ;
        RECT 22.300 84.240 37.630 84.470 ;
        RECT 15.720 83.325 16.450 83.355 ;
        RECT 15.720 83.255 16.510 83.325 ;
        RECT 15.700 82.835 16.510 83.255 ;
        RECT 15.720 82.785 16.510 82.835 ;
        RECT 15.720 82.755 16.450 82.785 ;
        RECT 18.820 81.955 19.760 82.545 ;
        RECT 17.500 80.695 18.320 80.725 ;
        RECT 15.270 80.615 15.620 80.665 ;
        RECT 15.010 80.585 15.620 80.615 ;
        RECT 14.980 80.415 15.640 80.585 ;
        RECT 14.980 79.985 15.620 80.415 ;
        RECT 17.500 80.225 18.340 80.695 ;
        RECT 17.500 80.195 18.320 80.225 ;
        RECT 15.000 79.945 15.620 79.985 ;
        RECT 17.790 79.715 18.130 80.195 ;
        RECT 17.780 79.555 18.130 79.715 ;
        RECT 17.770 79.475 18.130 79.555 ;
        RECT 17.770 79.285 18.120 79.475 ;
        RECT 17.770 79.165 18.170 79.285 ;
        RECT 17.800 79.045 18.170 79.165 ;
        RECT 17.800 78.985 18.150 79.045 ;
        RECT 23.000 73.830 23.230 84.240 ;
        RECT 23.440 74.030 23.710 84.040 ;
        RECT 25.020 74.030 25.290 84.040 ;
        RECT 26.600 74.030 26.870 84.040 ;
        RECT 28.180 74.030 28.450 84.040 ;
        RECT 29.760 74.030 30.030 84.040 ;
        RECT 31.340 74.030 31.610 84.040 ;
        RECT 32.920 74.030 33.190 84.040 ;
        RECT 34.500 74.030 34.770 84.040 ;
        RECT 36.080 74.030 36.350 84.040 ;
        RECT 37.660 74.030 37.930 84.040 ;
        RECT 121.200 83.800 121.430 85.210 ;
        RECT 106.100 83.570 121.430 83.800 ;
        RECT 23.000 73.600 37.630 73.830 ;
        RECT 105.800 73.360 106.070 83.370 ;
        RECT 107.380 73.360 107.650 83.370 ;
        RECT 108.960 73.360 109.230 83.370 ;
        RECT 110.540 73.360 110.810 83.370 ;
        RECT 112.120 73.360 112.390 83.370 ;
        RECT 113.700 73.360 113.970 83.370 ;
        RECT 115.280 73.360 115.550 83.370 ;
        RECT 116.860 73.360 117.130 83.370 ;
        RECT 118.440 73.360 118.710 83.370 ;
        RECT 120.020 73.360 120.290 83.370 ;
        RECT 120.500 73.160 120.730 83.570 ;
        RECT 127.280 82.655 128.010 82.685 ;
        RECT 127.220 82.585 128.010 82.655 ;
        RECT 127.220 82.165 128.030 82.585 ;
        RECT 127.220 82.115 128.010 82.165 ;
        RECT 127.280 82.085 128.010 82.115 ;
        RECT 123.970 81.285 124.910 81.875 ;
        RECT 125.410 80.025 126.230 80.055 ;
        RECT 125.390 79.555 126.230 80.025 ;
        RECT 128.110 79.945 128.460 79.995 ;
        RECT 128.110 79.915 128.720 79.945 ;
        RECT 128.090 79.745 128.750 79.915 ;
        RECT 125.410 79.525 126.230 79.555 ;
        RECT 125.600 79.045 125.940 79.525 ;
        RECT 128.110 79.315 128.750 79.745 ;
        RECT 128.110 79.275 128.730 79.315 ;
        RECT 125.600 78.885 125.950 79.045 ;
        RECT 125.600 78.805 125.960 78.885 ;
        RECT 125.610 78.615 125.960 78.805 ;
        RECT 125.560 78.495 125.960 78.615 ;
        RECT 125.560 78.375 125.930 78.495 ;
        RECT 125.580 78.315 125.930 78.375 ;
        RECT 106.100 72.930 120.730 73.160 ;
        RECT 23.255 66.465 37.885 66.695 ;
        RECT 22.955 56.255 23.225 66.265 ;
        RECT 24.535 56.255 24.805 66.265 ;
        RECT 26.115 56.255 26.385 66.265 ;
        RECT 27.695 56.255 27.965 66.265 ;
        RECT 29.275 56.255 29.545 66.265 ;
        RECT 30.855 56.255 31.125 66.265 ;
        RECT 32.435 56.255 32.705 66.265 ;
        RECT 34.015 56.255 34.285 66.265 ;
        RECT 35.595 56.255 35.865 66.265 ;
        RECT 37.175 56.255 37.445 66.265 ;
        RECT 37.655 56.055 37.885 66.465 ;
        RECT 104.855 66.465 119.485 66.695 ;
        RECT 104.855 56.055 105.085 66.465 ;
        RECT 105.295 56.255 105.565 66.265 ;
        RECT 106.875 56.255 107.145 66.265 ;
        RECT 108.455 56.255 108.725 66.265 ;
        RECT 110.035 56.255 110.305 66.265 ;
        RECT 111.615 56.255 111.885 66.265 ;
        RECT 113.195 56.255 113.465 66.265 ;
        RECT 114.775 56.255 115.045 66.265 ;
        RECT 116.355 56.255 116.625 66.265 ;
        RECT 117.935 56.255 118.205 66.265 ;
        RECT 119.515 56.255 119.785 66.265 ;
        RECT 23.255 55.825 38.585 56.055 ;
        RECT 38.355 54.415 38.585 55.825 ;
        RECT 35.045 54.185 38.585 54.415 ;
        RECT 104.155 55.825 119.485 56.055 ;
        RECT 104.155 54.415 104.385 55.825 ;
        RECT 104.155 54.185 107.695 54.415 ;
        RECT 23.105 52.895 32.995 53.125 ;
        RECT 22.805 47.735 23.075 52.735 ;
        RECT 24.385 47.735 24.655 52.735 ;
        RECT 25.965 47.735 26.235 52.735 ;
        RECT 27.545 47.735 27.815 52.735 ;
        RECT 29.125 47.735 29.395 52.735 ;
        RECT 30.705 47.735 30.975 52.735 ;
        RECT 32.285 47.735 32.555 52.735 ;
        RECT 32.765 50.115 32.995 52.895 ;
        RECT 35.045 52.905 35.275 54.185 ;
        RECT 37.875 53.695 39.165 53.925 ;
        RECT 36.145 52.905 36.375 53.575 ;
        RECT 35.045 52.655 36.375 52.905 ;
        RECT 37.825 52.665 38.795 52.895 ;
        RECT 36.145 51.985 36.375 52.655 ;
        RECT 37.525 51.585 38.415 51.815 ;
        RECT 36.145 50.115 36.375 50.785 ;
        RECT 32.765 49.865 36.375 50.115 ;
        RECT 37.525 50.105 37.755 51.585 ;
        RECT 38.555 51.185 38.795 52.665 ;
        RECT 37.895 50.955 38.795 51.185 ;
        RECT 37.525 49.875 38.485 50.105 ;
        RECT 32.765 47.575 32.995 49.865 ;
        RECT 36.145 49.195 36.375 49.865 ;
        RECT 37.875 48.845 38.525 49.075 ;
        RECT 37.875 48.615 38.045 48.845 ;
        RECT 23.105 47.345 32.995 47.575 ;
        RECT 36.635 48.445 38.045 48.615 ;
        RECT 34.645 46.495 34.965 46.555 ;
        RECT 36.635 46.495 36.805 48.445 ;
        RECT 38.995 47.835 39.165 53.695 ;
        RECT 37.015 47.545 39.165 47.835 ;
        RECT 103.575 53.695 104.865 53.925 ;
        RECT 103.575 47.835 103.745 53.695 ;
        RECT 106.365 52.905 106.595 53.575 ;
        RECT 107.465 52.905 107.695 54.185 ;
        RECT 103.945 52.665 104.915 52.895 ;
        RECT 103.945 51.185 104.185 52.665 ;
        RECT 106.365 52.655 107.695 52.905 ;
        RECT 109.745 52.895 119.635 53.125 ;
        RECT 106.365 51.985 106.595 52.655 ;
        RECT 104.325 51.585 105.215 51.815 ;
        RECT 103.945 50.955 104.845 51.185 ;
        RECT 104.985 50.105 105.215 51.585 ;
        RECT 104.255 49.875 105.215 50.105 ;
        RECT 106.365 50.115 106.595 50.785 ;
        RECT 109.745 50.115 109.975 52.895 ;
        RECT 106.365 49.865 109.975 50.115 ;
        RECT 106.365 49.195 106.595 49.865 ;
        RECT 104.215 48.845 104.865 49.075 ;
        RECT 104.695 48.615 104.865 48.845 ;
        RECT 104.695 48.445 106.105 48.615 ;
        RECT 103.575 47.545 105.725 47.835 ;
        RECT 37.595 47.115 37.825 47.405 ;
        RECT 104.915 47.115 105.145 47.405 ;
        RECT 37.625 46.495 37.795 47.115 ;
        RECT 34.645 46.325 37.795 46.495 ;
        RECT 104.945 46.495 105.115 47.115 ;
        RECT 105.935 46.495 106.105 48.445 ;
        RECT 109.745 47.575 109.975 49.865 ;
        RECT 110.185 47.735 110.455 52.735 ;
        RECT 111.765 47.735 112.035 52.735 ;
        RECT 113.345 47.735 113.615 52.735 ;
        RECT 114.925 47.735 115.195 52.735 ;
        RECT 116.505 47.735 116.775 52.735 ;
        RECT 118.085 47.735 118.355 52.735 ;
        RECT 119.665 47.735 119.935 52.735 ;
        RECT 109.745 47.345 119.635 47.575 ;
        RECT 107.775 46.495 108.095 46.555 ;
        RECT 104.945 46.325 108.095 46.495 ;
        RECT 34.645 46.295 34.965 46.325 ;
        RECT 107.775 46.295 108.095 46.325 ;
        RECT 99.380 44.575 102.250 44.690 ;
        RECT 39.920 44.555 41.290 44.575 ;
        RECT 39.920 44.550 41.460 44.555 ;
        RECT 39.920 44.545 45.630 44.550 ;
        RECT 38.930 43.480 45.630 44.545 ;
        RECT 99.380 44.545 102.820 44.575 ;
        RECT 99.380 44.530 103.810 44.545 ;
        RECT 38.930 43.475 41.290 43.480 ;
        RECT 38.930 43.445 40.300 43.475 ;
        RECT 18.660 43.405 19.320 43.425 ;
        RECT 19.520 43.405 21.440 43.425 ;
        RECT 18.660 43.400 22.830 43.405 ;
        RECT 25.590 43.400 25.910 43.430 ;
        RECT 18.660 43.230 25.910 43.400 ;
        RECT 18.660 43.215 22.930 43.230 ;
        RECT 18.660 42.815 19.320 43.215 ;
        RECT 19.520 43.205 21.440 43.215 ;
        RECT 22.760 42.610 22.930 43.215 ;
        RECT 22.730 42.320 22.960 42.610 ;
        RECT 21.390 41.890 23.540 42.180 ;
        RECT 13.910 37.365 14.570 38.385 ;
        RECT 18.850 37.925 19.640 38.625 ;
        RECT 13.970 35.335 14.610 36.355 ;
        RECT 21.390 36.030 21.560 41.890 ;
        RECT 23.750 41.280 23.920 43.230 ;
        RECT 25.590 43.170 25.910 43.230 ;
        RECT 22.510 41.110 23.920 41.280 ;
        RECT 27.560 42.150 37.450 42.380 ;
        RECT 22.510 40.880 22.680 41.110 ;
        RECT 22.030 40.650 22.680 40.880 ;
        RECT 24.180 39.860 24.410 40.530 ;
        RECT 27.560 39.860 27.790 42.150 ;
        RECT 22.070 39.620 23.030 39.850 ;
        RECT 21.760 38.540 22.660 38.770 ;
        RECT 21.760 37.060 22.000 38.540 ;
        RECT 22.800 38.140 23.030 39.620 ;
        RECT 24.180 39.610 27.790 39.860 ;
        RECT 24.180 38.940 24.410 39.610 ;
        RECT 22.140 37.910 23.030 38.140 ;
        RECT 24.180 37.070 24.410 37.740 ;
        RECT 21.760 36.830 22.730 37.060 ;
        RECT 24.180 36.820 25.510 37.070 ;
        RECT 24.180 36.150 24.410 36.820 ;
        RECT 21.390 35.800 22.680 36.030 ;
        RECT 25.280 35.540 25.510 36.820 ;
        RECT 27.560 36.830 27.790 39.610 ;
        RECT 28.000 36.990 28.270 41.990 ;
        RECT 29.580 36.990 29.850 41.990 ;
        RECT 31.160 36.990 31.430 41.990 ;
        RECT 32.740 36.990 33.010 41.990 ;
        RECT 34.320 36.990 34.590 41.990 ;
        RECT 35.900 36.990 36.170 41.990 ;
        RECT 37.480 36.990 37.750 41.990 ;
        RECT 27.560 36.600 37.450 36.830 ;
        RECT 42.880 35.650 44.920 43.480 ;
        RECT 96.450 43.475 103.810 44.530 ;
        RECT 96.450 43.460 102.250 43.475 ;
        RECT 97.160 35.630 99.200 43.460 ;
        RECT 99.380 43.410 102.250 43.460 ;
        RECT 102.440 43.445 103.810 43.475 ;
        RECT 116.830 43.400 117.150 43.430 ;
        RECT 121.300 43.405 123.220 43.425 ;
        RECT 123.420 43.405 124.080 43.425 ;
        RECT 119.910 43.400 124.080 43.405 ;
        RECT 116.830 43.230 124.080 43.400 ;
        RECT 116.830 43.170 117.150 43.230 ;
        RECT 105.290 42.150 115.180 42.380 ;
        RECT 104.990 36.990 105.260 41.990 ;
        RECT 106.570 36.990 106.840 41.990 ;
        RECT 108.150 36.990 108.420 41.990 ;
        RECT 109.730 36.990 110.000 41.990 ;
        RECT 111.310 36.990 111.580 41.990 ;
        RECT 112.890 36.990 113.160 41.990 ;
        RECT 114.470 36.990 114.740 41.990 ;
        RECT 114.950 39.860 115.180 42.150 ;
        RECT 118.820 41.280 118.990 43.230 ;
        RECT 119.810 43.215 124.080 43.230 ;
        RECT 119.810 42.610 119.980 43.215 ;
        RECT 121.300 43.205 123.220 43.215 ;
        RECT 123.420 42.815 124.080 43.215 ;
        RECT 119.780 42.320 120.010 42.610 ;
        RECT 119.200 41.890 121.350 42.180 ;
        RECT 118.820 41.110 120.230 41.280 ;
        RECT 120.060 40.880 120.230 41.110 ;
        RECT 120.060 40.650 120.710 40.880 ;
        RECT 118.330 39.860 118.560 40.530 ;
        RECT 114.950 39.610 118.560 39.860 ;
        RECT 114.950 36.830 115.180 39.610 ;
        RECT 118.330 38.940 118.560 39.610 ;
        RECT 119.710 39.620 120.670 39.850 ;
        RECT 119.710 38.140 119.940 39.620 ;
        RECT 120.080 38.540 120.980 38.770 ;
        RECT 119.710 37.910 120.600 38.140 ;
        RECT 118.330 37.070 118.560 37.740 ;
        RECT 105.290 36.600 115.180 36.830 ;
        RECT 117.230 36.820 118.560 37.070 ;
        RECT 120.740 37.060 120.980 38.540 ;
        RECT 120.010 36.830 120.980 37.060 ;
        RECT 21.970 35.310 25.510 35.540 ;
        RECT 117.230 35.540 117.460 36.820 ;
        RECT 118.330 36.150 118.560 36.820 ;
        RECT 121.180 36.030 121.350 41.890 ;
        RECT 123.100 37.925 123.890 38.625 ;
        RECT 128.170 37.365 128.830 38.385 ;
        RECT 120.060 35.800 121.350 36.030 ;
        RECT 117.230 35.310 120.770 35.540 ;
        RECT 128.130 35.335 128.770 36.355 ;
        RECT 21.970 33.900 22.200 35.310 ;
        RECT 120.540 33.900 120.770 35.310 ;
        RECT 21.970 33.670 37.300 33.900 ;
        RECT 105.440 33.670 120.770 33.900 ;
        RECT 15.390 32.755 16.120 32.785 ;
        RECT 15.390 32.685 16.180 32.755 ;
        RECT 15.370 32.265 16.180 32.685 ;
        RECT 15.390 32.215 16.180 32.265 ;
        RECT 15.390 32.185 16.120 32.215 ;
        RECT 18.490 31.385 19.430 31.975 ;
        RECT 17.170 30.125 17.990 30.155 ;
        RECT 14.940 30.045 15.290 30.095 ;
        RECT 14.680 30.015 15.290 30.045 ;
        RECT 14.650 29.845 15.310 30.015 ;
        RECT 14.650 29.415 15.290 29.845 ;
        RECT 17.170 29.655 18.010 30.125 ;
        RECT 17.170 29.625 17.990 29.655 ;
        RECT 14.670 29.375 15.290 29.415 ;
        RECT 17.460 29.145 17.800 29.625 ;
        RECT 17.450 28.985 17.800 29.145 ;
        RECT 17.440 28.905 17.800 28.985 ;
        RECT 17.440 28.715 17.790 28.905 ;
        RECT 17.440 28.595 17.840 28.715 ;
        RECT 17.470 28.475 17.840 28.595 ;
        RECT 17.470 28.415 17.820 28.475 ;
        RECT 22.670 23.260 22.900 33.670 ;
        RECT 23.110 23.460 23.380 33.470 ;
        RECT 24.690 23.460 24.960 33.470 ;
        RECT 26.270 23.460 26.540 33.470 ;
        RECT 27.850 23.460 28.120 33.470 ;
        RECT 29.430 23.460 29.700 33.470 ;
        RECT 31.010 23.460 31.280 33.470 ;
        RECT 32.590 23.460 32.860 33.470 ;
        RECT 34.170 23.460 34.440 33.470 ;
        RECT 35.750 23.460 36.020 33.470 ;
        RECT 37.330 23.460 37.600 33.470 ;
        RECT 105.140 23.460 105.410 33.470 ;
        RECT 106.720 23.460 106.990 33.470 ;
        RECT 108.300 23.460 108.570 33.470 ;
        RECT 109.880 23.460 110.150 33.470 ;
        RECT 111.460 23.460 111.730 33.470 ;
        RECT 113.040 23.460 113.310 33.470 ;
        RECT 114.620 23.460 114.890 33.470 ;
        RECT 116.200 23.460 116.470 33.470 ;
        RECT 117.780 23.460 118.050 33.470 ;
        RECT 119.360 23.460 119.630 33.470 ;
        RECT 119.840 23.260 120.070 33.670 ;
        RECT 126.620 32.755 127.350 32.785 ;
        RECT 126.560 32.685 127.350 32.755 ;
        RECT 126.560 32.265 127.370 32.685 ;
        RECT 126.560 32.215 127.350 32.265 ;
        RECT 126.620 32.185 127.350 32.215 ;
        RECT 123.310 31.385 124.250 31.975 ;
        RECT 124.750 30.125 125.570 30.155 ;
        RECT 124.730 29.655 125.570 30.125 ;
        RECT 127.450 30.045 127.800 30.095 ;
        RECT 127.450 30.015 128.060 30.045 ;
        RECT 127.430 29.845 128.090 30.015 ;
        RECT 124.750 29.625 125.570 29.655 ;
        RECT 124.940 29.145 125.280 29.625 ;
        RECT 127.450 29.415 128.090 29.845 ;
        RECT 127.450 29.375 128.070 29.415 ;
        RECT 124.940 28.985 125.290 29.145 ;
        RECT 124.940 28.905 125.300 28.985 ;
        RECT 124.950 28.715 125.300 28.905 ;
        RECT 124.900 28.595 125.300 28.715 ;
        RECT 124.900 28.475 125.270 28.595 ;
        RECT 124.920 28.415 125.270 28.475 ;
        RECT 22.670 23.030 37.300 23.260 ;
        RECT 105.440 23.030 120.070 23.260 ;
      LAYER met2 ;
        RECT 21.015 212.635 37.115 214.635 ;
        RECT 105.955 212.635 122.055 214.635 ;
        RECT 21.015 209.295 23.015 212.635 ;
        RECT 120.055 209.295 122.055 212.635 ;
        RECT 21.015 207.295 37.115 209.295 ;
        RECT 105.955 207.295 122.055 209.295 ;
        RECT 21.015 204.625 23.015 207.295 ;
        RECT 120.055 204.625 122.055 207.295 ;
        RECT 22.475 196.105 32.225 198.105 ;
        RECT 40.260 196.655 41.080 197.125 ;
        RECT 101.990 196.655 102.810 197.125 ;
        RECT 40.270 196.355 41.070 196.655 ;
        RECT 102.000 196.355 102.800 196.655 ;
        RECT 34.285 194.655 34.665 194.935 ;
        RECT 38.600 191.815 39.970 192.915 ;
        RECT 18.330 191.185 18.990 191.795 ;
        RECT 25.230 191.530 25.610 191.810 ;
        RECT 38.620 191.265 39.420 191.285 ;
        RECT 40.270 191.265 41.060 196.355 ;
        RECT 102.010 191.265 102.800 196.355 ;
        RECT 110.845 196.105 120.595 198.105 ;
        RECT 108.405 194.655 108.785 194.935 ;
        RECT 103.100 191.815 104.470 192.915 ;
        RECT 117.460 191.530 117.840 191.810 ;
        RECT 103.650 191.265 104.450 191.285 ;
        RECT 18.510 186.905 19.260 188.485 ;
        RECT 27.670 188.360 37.420 190.360 ;
        RECT 38.620 190.075 41.080 191.265 ;
        RECT 101.990 190.075 104.450 191.265 ;
        RECT 124.080 191.185 124.740 191.795 ;
        RECT 13.780 186.545 14.140 186.605 ;
        RECT 13.780 185.885 14.950 186.545 ;
        RECT 18.550 186.245 19.260 186.905 ;
        RECT 13.780 185.845 14.890 185.885 ;
        RECT 13.780 185.805 14.140 185.845 ;
        RECT 14.350 185.695 14.890 185.845 ;
        RECT 13.700 183.925 14.240 184.475 ;
        RECT 13.710 178.445 14.240 183.925 ;
        RECT 14.400 181.045 14.890 185.695 ;
        RECT 19.240 183.935 21.140 183.945 ;
        RECT 18.470 183.915 26.350 183.935 ;
        RECT 38.620 183.915 39.420 190.075 ;
        RECT 40.270 190.055 41.060 190.075 ;
        RECT 102.010 190.055 102.800 190.075 ;
        RECT 42.660 186.310 45.700 186.440 ;
        RECT 97.390 186.350 100.430 186.480 ;
        RECT 18.420 183.905 26.350 183.915 ;
        RECT 37.150 183.905 39.420 183.915 ;
        RECT 18.420 183.475 39.420 183.905 ;
        RECT 18.420 183.435 26.300 183.475 ;
        RECT 37.150 183.465 39.420 183.475 ;
        RECT 18.420 181.315 18.840 183.435 ;
        RECT 19.240 183.425 21.140 183.435 ;
        RECT 42.430 182.970 45.930 186.310 ;
        RECT 97.160 183.010 100.660 186.350 ;
        RECT 103.650 183.915 104.450 190.075 ;
        RECT 105.650 188.360 115.400 190.360 ;
        RECT 123.810 186.905 124.560 188.485 ;
        RECT 123.810 186.245 124.520 186.905 ;
        RECT 128.930 186.545 129.290 186.605 ;
        RECT 128.120 185.885 129.290 186.545 ;
        RECT 128.180 185.845 129.290 185.885 ;
        RECT 128.180 185.695 128.720 185.845 ;
        RECT 128.930 185.805 129.290 185.845 ;
        RECT 121.930 183.935 123.830 183.945 ;
        RECT 116.720 183.915 124.600 183.935 ;
        RECT 103.650 183.905 105.920 183.915 ;
        RECT 116.720 183.905 124.650 183.915 ;
        RECT 103.650 183.475 124.650 183.905 ;
        RECT 103.650 183.465 105.920 183.475 ;
        RECT 116.770 183.435 124.650 183.475 ;
        RECT 121.930 183.425 123.830 183.435 ;
        RECT 18.350 181.185 18.840 181.315 ;
        RECT 15.090 181.045 15.800 181.105 ;
        RECT 14.400 180.625 15.800 181.045 ;
        RECT 14.400 180.605 14.890 180.625 ;
        RECT 15.090 180.585 15.800 180.625 ;
        RECT 18.350 180.295 18.780 181.185 ;
        RECT 18.290 179.915 18.920 180.295 ;
        RECT 18.280 179.845 18.920 179.915 ;
        RECT 18.270 178.595 18.920 179.845 ;
        RECT 36.880 179.170 38.880 181.840 ;
        RECT 13.710 178.435 14.400 178.445 ;
        RECT 13.710 177.735 14.930 178.435 ;
        RECT 16.880 178.265 18.920 178.595 ;
        RECT 16.880 178.005 17.630 178.265 ;
        RECT 18.330 178.245 18.920 178.265 ;
        RECT 16.890 177.975 17.630 178.005 ;
        RECT 13.710 177.715 14.400 177.735 ;
        RECT 14.190 177.705 14.400 177.715 ;
        RECT 22.780 177.170 38.880 179.170 ;
        RECT 36.880 173.830 38.880 177.170 ;
        RECT 22.780 171.830 38.880 173.830 ;
        RECT 104.190 179.170 106.190 181.840 ;
        RECT 124.230 181.315 124.650 183.435 ;
        RECT 124.230 181.185 124.720 181.315 ;
        RECT 124.290 180.295 124.720 181.185 ;
        RECT 127.270 181.045 127.980 181.105 ;
        RECT 128.180 181.045 128.670 185.695 ;
        RECT 127.270 180.625 128.670 181.045 ;
        RECT 127.270 180.585 127.980 180.625 ;
        RECT 128.180 180.605 128.670 180.625 ;
        RECT 128.830 183.925 129.370 184.475 ;
        RECT 124.150 179.915 124.780 180.295 ;
        RECT 124.150 179.845 124.790 179.915 ;
        RECT 104.190 177.170 120.290 179.170 ;
        RECT 124.150 178.595 124.800 179.845 ;
        RECT 124.150 178.265 126.190 178.595 ;
        RECT 128.830 178.445 129.360 183.925 ;
        RECT 128.670 178.435 129.360 178.445 ;
        RECT 124.150 178.245 124.740 178.265 ;
        RECT 125.440 178.005 126.190 178.265 ;
        RECT 125.440 177.975 126.180 178.005 ;
        RECT 128.140 177.735 129.360 178.435 ;
        RECT 128.670 177.715 129.360 177.735 ;
        RECT 128.670 177.705 128.880 177.715 ;
        RECT 104.190 173.830 106.190 177.170 ;
        RECT 104.190 171.830 120.290 173.830 ;
        RECT 21.015 163.065 37.115 165.065 ;
        RECT 105.955 163.065 122.055 165.065 ;
        RECT 21.015 159.725 23.015 163.065 ;
        RECT 120.055 159.725 122.055 163.065 ;
        RECT 21.015 157.725 37.115 159.725 ;
        RECT 105.955 157.725 122.055 159.725 ;
        RECT 21.015 155.055 23.015 157.725 ;
        RECT 120.055 155.055 122.055 157.725 ;
        RECT 22.475 146.535 32.225 148.535 ;
        RECT 40.260 147.085 41.080 147.555 ;
        RECT 101.990 147.085 102.810 147.555 ;
        RECT 40.270 146.785 41.070 147.085 ;
        RECT 102.000 146.785 102.800 147.085 ;
        RECT 34.285 145.085 34.665 145.365 ;
        RECT 38.600 142.245 39.970 143.345 ;
        RECT 18.330 141.615 18.990 142.225 ;
        RECT 25.230 141.960 25.610 142.240 ;
        RECT 38.620 141.695 39.420 141.715 ;
        RECT 40.270 141.695 41.060 146.785 ;
        RECT 102.010 141.695 102.800 146.785 ;
        RECT 110.845 146.535 120.595 148.535 ;
        RECT 108.405 145.085 108.785 145.365 ;
        RECT 103.100 142.245 104.470 143.345 ;
        RECT 117.460 141.960 117.840 142.240 ;
        RECT 103.650 141.695 104.450 141.715 ;
        RECT 18.510 137.335 19.260 138.915 ;
        RECT 27.670 138.790 37.420 140.790 ;
        RECT 38.620 140.505 41.080 141.695 ;
        RECT 101.990 140.505 104.450 141.695 ;
        RECT 124.080 141.615 124.740 142.225 ;
        RECT 13.780 136.975 14.140 137.035 ;
        RECT 13.780 136.315 14.950 136.975 ;
        RECT 18.550 136.675 19.260 137.335 ;
        RECT 13.780 136.275 14.890 136.315 ;
        RECT 13.780 136.235 14.140 136.275 ;
        RECT 14.350 136.125 14.890 136.275 ;
        RECT 13.700 134.355 14.240 134.905 ;
        RECT 13.710 128.875 14.240 134.355 ;
        RECT 14.400 131.475 14.890 136.125 ;
        RECT 19.240 134.365 21.140 134.375 ;
        RECT 18.470 134.345 26.350 134.365 ;
        RECT 38.620 134.345 39.420 140.505 ;
        RECT 40.270 140.485 41.060 140.505 ;
        RECT 102.010 140.485 102.800 140.505 ;
        RECT 42.710 136.780 45.750 136.910 ;
        RECT 18.420 134.335 26.350 134.345 ;
        RECT 37.150 134.335 39.420 134.345 ;
        RECT 18.420 133.905 39.420 134.335 ;
        RECT 18.420 133.865 26.300 133.905 ;
        RECT 37.150 133.895 39.420 133.905 ;
        RECT 18.420 131.745 18.840 133.865 ;
        RECT 19.240 133.855 21.140 133.865 ;
        RECT 42.480 133.440 45.980 136.780 ;
        RECT 97.260 136.740 100.300 136.870 ;
        RECT 97.030 133.400 100.530 136.740 ;
        RECT 103.650 134.345 104.450 140.505 ;
        RECT 105.650 138.790 115.400 140.790 ;
        RECT 123.810 137.335 124.560 138.915 ;
        RECT 123.810 136.675 124.520 137.335 ;
        RECT 128.930 136.975 129.290 137.035 ;
        RECT 128.120 136.315 129.290 136.975 ;
        RECT 128.180 136.275 129.290 136.315 ;
        RECT 128.180 136.125 128.720 136.275 ;
        RECT 128.930 136.235 129.290 136.275 ;
        RECT 121.930 134.365 123.830 134.375 ;
        RECT 116.720 134.345 124.600 134.365 ;
        RECT 103.650 134.335 105.920 134.345 ;
        RECT 116.720 134.335 124.650 134.345 ;
        RECT 103.650 133.905 124.650 134.335 ;
        RECT 103.650 133.895 105.920 133.905 ;
        RECT 116.770 133.865 124.650 133.905 ;
        RECT 121.930 133.855 123.830 133.865 ;
        RECT 18.350 131.615 18.840 131.745 ;
        RECT 15.090 131.475 15.800 131.535 ;
        RECT 14.400 131.055 15.800 131.475 ;
        RECT 14.400 131.035 14.890 131.055 ;
        RECT 15.090 131.015 15.800 131.055 ;
        RECT 18.350 130.725 18.780 131.615 ;
        RECT 18.290 130.345 18.920 130.725 ;
        RECT 18.280 130.275 18.920 130.345 ;
        RECT 18.270 129.025 18.920 130.275 ;
        RECT 36.880 129.600 38.880 132.270 ;
        RECT 13.710 128.865 14.400 128.875 ;
        RECT 13.710 128.165 14.930 128.865 ;
        RECT 16.880 128.695 18.920 129.025 ;
        RECT 16.880 128.435 17.630 128.695 ;
        RECT 18.330 128.675 18.920 128.695 ;
        RECT 16.890 128.405 17.630 128.435 ;
        RECT 13.710 128.145 14.400 128.165 ;
        RECT 14.190 128.135 14.400 128.145 ;
        RECT 22.780 127.600 38.880 129.600 ;
        RECT 36.880 124.260 38.880 127.600 ;
        RECT 22.780 122.260 38.880 124.260 ;
        RECT 104.190 129.600 106.190 132.270 ;
        RECT 124.230 131.745 124.650 133.865 ;
        RECT 124.230 131.615 124.720 131.745 ;
        RECT 124.290 130.725 124.720 131.615 ;
        RECT 127.270 131.475 127.980 131.535 ;
        RECT 128.180 131.475 128.670 136.125 ;
        RECT 127.270 131.055 128.670 131.475 ;
        RECT 127.270 131.015 127.980 131.055 ;
        RECT 128.180 131.035 128.670 131.055 ;
        RECT 128.830 134.355 129.370 134.905 ;
        RECT 124.150 130.345 124.780 130.725 ;
        RECT 124.150 130.275 124.790 130.345 ;
        RECT 104.190 127.600 120.290 129.600 ;
        RECT 124.150 129.025 124.800 130.275 ;
        RECT 124.150 128.695 126.190 129.025 ;
        RECT 128.830 128.875 129.360 134.355 ;
        RECT 128.670 128.865 129.360 128.875 ;
        RECT 124.150 128.675 124.740 128.695 ;
        RECT 125.440 128.435 126.190 128.695 ;
        RECT 125.440 128.405 126.180 128.435 ;
        RECT 128.140 128.165 129.360 128.865 ;
        RECT 128.670 128.145 129.360 128.165 ;
        RECT 128.670 128.135 128.880 128.145 ;
        RECT 104.190 124.260 106.190 127.600 ;
        RECT 104.190 122.260 120.290 124.260 ;
        RECT 21.675 114.835 37.775 116.835 ;
        RECT 21.675 111.495 23.675 114.835 ;
        RECT 105.955 114.165 122.055 116.165 ;
        RECT 21.675 109.495 37.775 111.495 ;
        RECT 120.055 110.825 122.055 114.165 ;
        RECT 21.675 106.825 23.675 109.495 ;
        RECT 105.955 108.825 122.055 110.825 ;
        RECT 120.055 106.155 122.055 108.825 ;
        RECT 23.135 98.305 32.885 100.305 ;
        RECT 40.920 98.855 41.740 99.325 ;
        RECT 40.930 98.555 41.730 98.855 ;
        RECT 34.945 96.855 35.325 97.135 ;
        RECT 39.260 94.015 40.630 95.115 ;
        RECT 18.990 93.385 19.650 93.995 ;
        RECT 25.890 93.730 26.270 94.010 ;
        RECT 39.280 93.465 40.080 93.485 ;
        RECT 40.930 93.465 41.720 98.555 ;
        RECT 101.990 98.185 102.810 98.655 ;
        RECT 102.000 97.885 102.800 98.185 ;
        RECT 19.170 89.105 19.920 90.685 ;
        RECT 28.330 90.560 38.080 92.560 ;
        RECT 39.280 92.275 41.740 93.465 ;
        RECT 102.010 92.795 102.800 97.885 ;
        RECT 110.845 97.635 120.595 99.635 ;
        RECT 108.405 96.185 108.785 96.465 ;
        RECT 103.100 93.345 104.470 94.445 ;
        RECT 117.460 93.060 117.840 93.340 ;
        RECT 103.650 92.795 104.450 92.815 ;
        RECT 14.440 88.745 14.800 88.805 ;
        RECT 14.440 88.085 15.610 88.745 ;
        RECT 19.210 88.445 19.920 89.105 ;
        RECT 14.440 88.045 15.550 88.085 ;
        RECT 14.440 88.005 14.800 88.045 ;
        RECT 15.010 87.895 15.550 88.045 ;
        RECT 14.360 86.125 14.900 86.675 ;
        RECT 14.370 80.645 14.900 86.125 ;
        RECT 15.060 83.245 15.550 87.895 ;
        RECT 19.900 86.135 21.800 86.145 ;
        RECT 19.130 86.115 27.010 86.135 ;
        RECT 39.280 86.115 40.080 92.275 ;
        RECT 40.930 92.255 41.720 92.275 ;
        RECT 101.990 91.605 104.450 92.795 ;
        RECT 124.080 92.715 124.740 93.325 ;
        RECT 102.010 91.585 102.800 91.605 ;
        RECT 43.210 88.590 46.250 88.720 ;
        RECT 19.080 86.105 27.010 86.115 ;
        RECT 37.810 86.105 40.080 86.115 ;
        RECT 19.080 85.675 40.080 86.105 ;
        RECT 19.080 85.635 26.960 85.675 ;
        RECT 37.810 85.665 40.080 85.675 ;
        RECT 19.080 83.515 19.500 85.635 ;
        RECT 19.900 85.625 21.800 85.635 ;
        RECT 42.980 85.250 46.480 88.590 ;
        RECT 97.350 87.800 100.390 87.930 ;
        RECT 97.120 84.460 100.620 87.800 ;
        RECT 103.650 85.445 104.450 91.605 ;
        RECT 105.650 89.890 115.400 91.890 ;
        RECT 123.810 88.435 124.560 90.015 ;
        RECT 123.810 87.775 124.520 88.435 ;
        RECT 128.930 88.075 129.290 88.135 ;
        RECT 128.120 87.415 129.290 88.075 ;
        RECT 128.180 87.375 129.290 87.415 ;
        RECT 128.180 87.225 128.720 87.375 ;
        RECT 128.930 87.335 129.290 87.375 ;
        RECT 121.930 85.465 123.830 85.475 ;
        RECT 116.720 85.445 124.600 85.465 ;
        RECT 103.650 85.435 105.920 85.445 ;
        RECT 116.720 85.435 124.650 85.445 ;
        RECT 103.650 85.005 124.650 85.435 ;
        RECT 103.650 84.995 105.920 85.005 ;
        RECT 116.770 84.965 124.650 85.005 ;
        RECT 121.930 84.955 123.830 84.965 ;
        RECT 19.010 83.385 19.500 83.515 ;
        RECT 15.750 83.245 16.460 83.305 ;
        RECT 15.060 82.825 16.460 83.245 ;
        RECT 15.060 82.805 15.550 82.825 ;
        RECT 15.750 82.785 16.460 82.825 ;
        RECT 19.010 82.495 19.440 83.385 ;
        RECT 18.950 82.115 19.580 82.495 ;
        RECT 18.940 82.045 19.580 82.115 ;
        RECT 18.930 80.795 19.580 82.045 ;
        RECT 37.540 81.370 39.540 84.040 ;
        RECT 14.370 80.635 15.060 80.645 ;
        RECT 14.370 79.935 15.590 80.635 ;
        RECT 17.540 80.465 19.580 80.795 ;
        RECT 17.540 80.205 18.290 80.465 ;
        RECT 18.990 80.445 19.580 80.465 ;
        RECT 17.550 80.175 18.290 80.205 ;
        RECT 14.370 79.915 15.060 79.935 ;
        RECT 14.850 79.905 15.060 79.915 ;
        RECT 23.440 79.370 39.540 81.370 ;
        RECT 37.540 76.030 39.540 79.370 ;
        RECT 23.440 74.030 39.540 76.030 ;
        RECT 104.190 80.700 106.190 83.370 ;
        RECT 124.230 82.845 124.650 84.965 ;
        RECT 124.230 82.715 124.720 82.845 ;
        RECT 124.290 81.825 124.720 82.715 ;
        RECT 127.270 82.575 127.980 82.635 ;
        RECT 128.180 82.575 128.670 87.225 ;
        RECT 127.270 82.155 128.670 82.575 ;
        RECT 127.270 82.115 127.980 82.155 ;
        RECT 128.180 82.135 128.670 82.155 ;
        RECT 128.830 85.455 129.370 86.005 ;
        RECT 124.150 81.445 124.780 81.825 ;
        RECT 124.150 81.375 124.790 81.445 ;
        RECT 104.190 78.700 120.290 80.700 ;
        RECT 124.150 80.125 124.800 81.375 ;
        RECT 124.150 79.795 126.190 80.125 ;
        RECT 128.830 79.975 129.360 85.455 ;
        RECT 128.670 79.965 129.360 79.975 ;
        RECT 124.150 79.775 124.740 79.795 ;
        RECT 125.440 79.535 126.190 79.795 ;
        RECT 125.440 79.505 126.180 79.535 ;
        RECT 128.140 79.265 129.360 79.965 ;
        RECT 128.670 79.245 129.360 79.265 ;
        RECT 128.670 79.235 128.880 79.245 ;
        RECT 104.190 75.360 106.190 78.700 ;
        RECT 104.190 73.360 120.290 75.360 ;
        RECT 21.345 64.265 37.445 66.265 ;
        RECT 105.295 64.265 121.395 66.265 ;
        RECT 21.345 60.925 23.345 64.265 ;
        RECT 119.395 60.925 121.395 64.265 ;
        RECT 21.345 58.925 37.445 60.925 ;
        RECT 105.295 58.925 121.395 60.925 ;
        RECT 21.345 56.255 23.345 58.925 ;
        RECT 119.395 56.255 121.395 58.925 ;
        RECT 22.805 47.735 32.555 49.735 ;
        RECT 40.590 48.285 41.410 48.755 ;
        RECT 101.330 48.285 102.150 48.755 ;
        RECT 40.600 47.985 41.400 48.285 ;
        RECT 101.340 47.985 102.140 48.285 ;
        RECT 34.615 46.285 34.995 46.565 ;
        RECT 38.930 43.445 40.300 44.545 ;
        RECT 18.660 42.815 19.320 43.425 ;
        RECT 25.560 43.160 25.940 43.440 ;
        RECT 38.950 42.895 39.750 42.915 ;
        RECT 40.600 42.895 41.390 47.985 ;
        RECT 101.350 42.895 102.140 47.985 ;
        RECT 110.185 47.735 119.935 49.735 ;
        RECT 107.745 46.285 108.125 46.565 ;
        RECT 102.440 43.445 103.810 44.545 ;
        RECT 116.800 43.160 117.180 43.440 ;
        RECT 102.990 42.895 103.790 42.915 ;
        RECT 18.840 38.535 19.590 40.115 ;
        RECT 28.000 39.990 37.750 41.990 ;
        RECT 38.950 41.705 41.410 42.895 ;
        RECT 101.330 41.705 103.790 42.895 ;
        RECT 123.420 42.815 124.080 43.425 ;
        RECT 14.110 38.175 14.470 38.235 ;
        RECT 14.110 37.515 15.280 38.175 ;
        RECT 18.880 37.875 19.590 38.535 ;
        RECT 14.110 37.475 15.220 37.515 ;
        RECT 14.110 37.435 14.470 37.475 ;
        RECT 14.680 37.325 15.220 37.475 ;
        RECT 14.030 35.555 14.570 36.105 ;
        RECT 14.040 30.075 14.570 35.555 ;
        RECT 14.730 32.675 15.220 37.325 ;
        RECT 19.570 35.565 21.470 35.575 ;
        RECT 18.800 35.545 26.680 35.565 ;
        RECT 38.950 35.545 39.750 41.705 ;
        RECT 40.600 41.685 41.390 41.705 ;
        RECT 101.350 41.685 102.140 41.705 ;
        RECT 42.700 37.990 45.740 38.120 ;
        RECT 18.750 35.535 26.680 35.545 ;
        RECT 37.480 35.535 39.750 35.545 ;
        RECT 18.750 35.105 39.750 35.535 ;
        RECT 18.750 35.065 26.630 35.105 ;
        RECT 37.480 35.095 39.750 35.105 ;
        RECT 18.750 32.945 19.170 35.065 ;
        RECT 19.570 35.055 21.470 35.065 ;
        RECT 42.470 34.650 45.970 37.990 ;
        RECT 96.340 37.970 99.380 38.100 ;
        RECT 96.110 34.630 99.610 37.970 ;
        RECT 102.990 35.545 103.790 41.705 ;
        RECT 104.990 39.990 114.740 41.990 ;
        RECT 123.150 38.535 123.900 40.115 ;
        RECT 123.150 37.875 123.860 38.535 ;
        RECT 128.270 38.175 128.630 38.235 ;
        RECT 127.460 37.515 128.630 38.175 ;
        RECT 127.520 37.475 128.630 37.515 ;
        RECT 127.520 37.325 128.060 37.475 ;
        RECT 128.270 37.435 128.630 37.475 ;
        RECT 121.270 35.565 123.170 35.575 ;
        RECT 116.060 35.545 123.940 35.565 ;
        RECT 102.990 35.535 105.260 35.545 ;
        RECT 116.060 35.535 123.990 35.545 ;
        RECT 102.990 35.105 123.990 35.535 ;
        RECT 102.990 35.095 105.260 35.105 ;
        RECT 116.110 35.065 123.990 35.105 ;
        RECT 121.270 35.055 123.170 35.065 ;
        RECT 18.680 32.815 19.170 32.945 ;
        RECT 15.420 32.675 16.130 32.735 ;
        RECT 14.730 32.255 16.130 32.675 ;
        RECT 14.730 32.235 15.220 32.255 ;
        RECT 15.420 32.215 16.130 32.255 ;
        RECT 18.680 31.925 19.110 32.815 ;
        RECT 18.620 31.545 19.250 31.925 ;
        RECT 18.610 31.475 19.250 31.545 ;
        RECT 18.600 30.225 19.250 31.475 ;
        RECT 37.210 30.800 39.210 33.470 ;
        RECT 14.040 30.065 14.730 30.075 ;
        RECT 14.040 29.365 15.260 30.065 ;
        RECT 17.210 29.895 19.250 30.225 ;
        RECT 17.210 29.635 17.960 29.895 ;
        RECT 18.660 29.875 19.250 29.895 ;
        RECT 17.220 29.605 17.960 29.635 ;
        RECT 14.040 29.345 14.730 29.365 ;
        RECT 14.520 29.335 14.730 29.345 ;
        RECT 23.110 28.800 39.210 30.800 ;
        RECT 37.210 25.460 39.210 28.800 ;
        RECT 23.110 23.460 39.210 25.460 ;
        RECT 103.530 30.800 105.530 33.470 ;
        RECT 123.570 32.945 123.990 35.065 ;
        RECT 123.570 32.815 124.060 32.945 ;
        RECT 123.630 31.925 124.060 32.815 ;
        RECT 126.610 32.675 127.320 32.735 ;
        RECT 127.520 32.675 128.010 37.325 ;
        RECT 126.610 32.255 128.010 32.675 ;
        RECT 126.610 32.215 127.320 32.255 ;
        RECT 127.520 32.235 128.010 32.255 ;
        RECT 128.170 35.555 128.710 36.105 ;
        RECT 123.490 31.545 124.120 31.925 ;
        RECT 123.490 31.475 124.130 31.545 ;
        RECT 103.530 28.800 119.630 30.800 ;
        RECT 123.490 30.225 124.140 31.475 ;
        RECT 123.490 29.895 125.530 30.225 ;
        RECT 128.170 30.075 128.700 35.555 ;
        RECT 128.010 30.065 128.700 30.075 ;
        RECT 123.490 29.875 124.080 29.895 ;
        RECT 124.780 29.635 125.530 29.895 ;
        RECT 124.780 29.605 125.520 29.635 ;
        RECT 127.480 29.365 128.700 30.065 ;
        RECT 128.010 29.345 128.700 29.365 ;
        RECT 128.010 29.335 128.220 29.345 ;
        RECT 103.530 25.460 105.530 28.800 ;
        RECT 103.530 23.460 119.630 25.460 ;
      LAYER met3 ;
        RECT 62.540 210.000 73.540 210.080 ;
        RECT 21.015 198.105 23.015 207.295 ;
        RECT 62.540 203.620 84.430 210.000 ;
        RECT 58.620 203.580 95.350 203.620 ;
        RECT 58.540 199.580 95.350 203.580 ;
        RECT 62.540 199.500 95.350 199.580 ;
        RECT 62.540 199.080 84.430 199.500 ;
        RECT 73.430 199.000 84.430 199.080 ;
        RECT 120.055 198.105 122.055 207.295 ;
        RECT 21.015 196.105 32.225 198.105 ;
        RECT 34.880 196.975 35.870 197.045 ;
        RECT 40.320 197.035 41.000 197.070 ;
        RECT 38.190 196.985 41.000 197.035 ;
        RECT 34.610 196.865 35.870 196.975 ;
        RECT 37.680 196.865 41.000 196.985 ;
        RECT 34.610 196.515 41.000 196.865 ;
        RECT 34.610 196.495 37.890 196.515 ;
        RECT 40.320 196.500 41.000 196.515 ;
        RECT 34.610 195.505 34.910 196.495 ;
        RECT 34.325 194.985 34.910 195.505 ;
        RECT 34.305 194.935 34.910 194.985 ;
        RECT 34.305 194.605 34.645 194.935 ;
        RECT 18.340 191.785 18.860 191.795 ;
        RECT 18.340 191.185 19.010 191.785 ;
        RECT 25.250 191.480 25.590 191.860 ;
        RECT 38.600 191.815 39.970 192.915 ;
        RECT 38.600 191.765 39.910 191.815 ;
        RECT 18.600 191.035 19.010 191.185 ;
        RECT 18.600 190.825 19.020 191.035 ;
        RECT 25.270 190.960 25.570 191.480 ;
        RECT 17.570 190.785 19.020 190.825 ;
        RECT 17.550 190.565 19.020 190.785 ;
        RECT 17.550 190.505 19.010 190.565 ;
        RECT 17.550 190.435 17.990 190.505 ;
        RECT 17.550 188.865 17.980 190.435 ;
        RECT 17.550 188.545 19.160 188.865 ;
        RECT 17.560 188.355 19.160 188.545 ;
        RECT 27.670 188.360 38.880 190.360 ;
        RECT 18.550 187.915 19.160 188.355 ;
        RECT 18.570 187.790 19.150 187.915 ;
        RECT 36.880 179.170 38.880 188.360 ;
        RECT 41.740 186.330 52.740 197.330 ;
        RECT 90.350 186.370 101.350 197.370 ;
        RECT 102.070 197.035 102.750 197.070 ;
        RECT 102.070 196.985 104.880 197.035 ;
        RECT 102.070 196.865 105.390 196.985 ;
        RECT 107.200 196.975 108.190 197.045 ;
        RECT 107.200 196.865 108.460 196.975 ;
        RECT 102.070 196.515 108.460 196.865 ;
        RECT 102.070 196.500 102.750 196.515 ;
        RECT 105.180 196.495 108.460 196.515 ;
        RECT 108.160 195.505 108.460 196.495 ;
        RECT 110.845 196.105 122.055 198.105 ;
        RECT 108.160 194.985 108.745 195.505 ;
        RECT 108.160 194.935 108.765 194.985 ;
        RECT 108.425 194.605 108.765 194.935 ;
        RECT 103.100 191.815 104.470 192.915 ;
        RECT 103.160 191.765 104.470 191.815 ;
        RECT 117.480 191.480 117.820 191.860 ;
        RECT 124.210 191.785 124.730 191.795 ;
        RECT 117.500 190.960 117.800 191.480 ;
        RECT 124.060 191.185 124.730 191.785 ;
        RECT 124.060 191.035 124.470 191.185 ;
        RECT 124.050 190.825 124.470 191.035 ;
        RECT 124.050 190.785 125.500 190.825 ;
        RECT 124.050 190.565 125.520 190.785 ;
        RECT 124.060 190.505 125.520 190.565 ;
        RECT 125.080 190.435 125.520 190.505 ;
        RECT 104.190 188.360 115.400 190.360 ;
        RECT 125.090 188.865 125.520 190.435 ;
        RECT 123.910 188.545 125.520 188.865 ;
        RECT 42.240 182.330 46.240 186.330 ;
        RECT 52.660 179.840 61.280 183.960 ;
        RECT 96.850 182.370 100.850 186.370 ;
        RECT 97.170 180.910 101.150 180.930 ;
        RECT 52.660 176.170 56.780 179.840 ;
        RECT 97.170 176.910 101.290 180.910 ;
        RECT 104.190 179.170 106.190 188.360 ;
        RECT 123.910 188.355 125.510 188.545 ;
        RECT 123.910 187.915 124.520 188.355 ;
        RECT 123.920 187.790 124.500 187.915 ;
        RECT 46.280 165.280 57.280 176.170 ;
        RECT 90.790 166.020 101.790 176.910 ;
        RECT 46.200 165.170 57.280 165.280 ;
        RECT 90.710 165.910 101.790 166.020 ;
        RECT 21.015 148.535 23.015 157.725 ;
        RECT 46.200 154.280 57.200 165.170 ;
        RECT 90.710 155.140 101.710 165.910 ;
        RECT 84.270 155.020 101.710 155.140 ;
        RECT 52.660 150.360 56.700 154.280 ;
        RECT 52.700 150.280 56.700 150.360 ;
        RECT 84.270 151.100 101.210 155.020 ;
        RECT 21.015 146.535 32.225 148.535 ;
        RECT 34.880 147.405 35.870 147.475 ;
        RECT 40.320 147.465 41.000 147.500 ;
        RECT 38.190 147.415 41.000 147.465 ;
        RECT 34.610 147.295 35.870 147.405 ;
        RECT 37.680 147.295 41.000 147.415 ;
        RECT 34.610 146.945 41.000 147.295 ;
        RECT 34.610 146.925 37.890 146.945 ;
        RECT 40.320 146.930 41.000 146.945 ;
        RECT 34.610 145.935 34.910 146.925 ;
        RECT 34.325 145.415 34.910 145.935 ;
        RECT 34.305 145.365 34.910 145.415 ;
        RECT 34.305 145.035 34.645 145.365 ;
        RECT 18.340 142.215 18.860 142.225 ;
        RECT 18.340 141.615 19.010 142.215 ;
        RECT 25.250 141.910 25.590 142.290 ;
        RECT 38.600 142.245 39.970 143.345 ;
        RECT 38.600 142.195 39.910 142.245 ;
        RECT 18.600 141.465 19.010 141.615 ;
        RECT 18.600 141.255 19.020 141.465 ;
        RECT 25.270 141.390 25.570 141.910 ;
        RECT 17.570 141.215 19.020 141.255 ;
        RECT 17.550 140.995 19.020 141.215 ;
        RECT 17.550 140.935 19.010 140.995 ;
        RECT 17.550 140.865 17.990 140.935 ;
        RECT 17.550 139.295 17.980 140.865 ;
        RECT 17.550 138.975 19.160 139.295 ;
        RECT 17.560 138.785 19.160 138.975 ;
        RECT 27.670 138.790 38.880 140.790 ;
        RECT 18.550 138.345 19.160 138.785 ;
        RECT 18.570 138.220 19.150 138.345 ;
        RECT 36.880 129.600 38.880 138.790 ;
        RECT 41.790 136.800 52.790 147.800 ;
        RECT 84.270 138.040 88.310 151.100 ;
        RECT 97.210 151.020 101.210 151.100 ;
        RECT 120.055 148.535 122.055 157.725 ;
        RECT 42.290 132.800 46.290 136.800 ;
        RECT 90.220 136.760 101.220 147.760 ;
        RECT 102.070 147.465 102.750 147.500 ;
        RECT 102.070 147.415 104.880 147.465 ;
        RECT 102.070 147.295 105.390 147.415 ;
        RECT 107.200 147.405 108.190 147.475 ;
        RECT 107.200 147.295 108.460 147.405 ;
        RECT 102.070 146.945 108.460 147.295 ;
        RECT 102.070 146.930 102.750 146.945 ;
        RECT 105.180 146.925 108.460 146.945 ;
        RECT 108.160 145.935 108.460 146.925 ;
        RECT 110.845 146.535 122.055 148.535 ;
        RECT 108.160 145.415 108.745 145.935 ;
        RECT 108.160 145.365 108.765 145.415 ;
        RECT 108.425 145.035 108.765 145.365 ;
        RECT 103.100 142.245 104.470 143.345 ;
        RECT 103.160 142.195 104.470 142.245 ;
        RECT 117.480 141.910 117.820 142.290 ;
        RECT 124.210 142.215 124.730 142.225 ;
        RECT 117.500 141.390 117.800 141.910 ;
        RECT 124.060 141.615 124.730 142.215 ;
        RECT 124.060 141.465 124.470 141.615 ;
        RECT 124.050 141.255 124.470 141.465 ;
        RECT 124.050 141.215 125.500 141.255 ;
        RECT 124.050 140.995 125.520 141.215 ;
        RECT 124.060 140.935 125.520 140.995 ;
        RECT 125.080 140.865 125.520 140.935 ;
        RECT 104.190 138.790 115.400 140.790 ;
        RECT 125.090 139.295 125.520 140.865 ;
        RECT 123.910 138.975 125.520 139.295 ;
        RECT 96.720 132.760 100.720 136.760 ;
        RECT 52.250 131.780 56.250 131.830 ;
        RECT 52.210 127.830 56.250 131.780 ;
        RECT 96.720 130.780 100.720 130.860 ;
        RECT 45.750 116.940 56.750 127.830 ;
        RECT 96.680 126.860 100.720 130.780 ;
        RECT 104.190 129.600 106.190 138.790 ;
        RECT 123.910 138.785 125.510 138.975 ;
        RECT 123.910 138.345 124.520 138.785 ;
        RECT 123.920 138.220 124.500 138.345 ;
        RECT 45.750 116.830 56.830 116.940 ;
        RECT 21.675 100.305 23.675 109.495 ;
        RECT 45.830 105.940 56.830 116.830 ;
        RECT 90.220 115.970 101.220 126.860 ;
        RECT 90.220 115.860 101.300 115.970 ;
        RECT 52.210 101.940 56.330 105.940 ;
        RECT 83.460 105.090 87.580 105.120 ;
        RECT 90.300 105.090 101.300 115.860 ;
        RECT 83.460 104.970 101.300 105.090 ;
        RECT 52.210 101.920 56.190 101.940 ;
        RECT 83.460 100.970 100.800 104.970 ;
        RECT 83.460 100.940 87.580 100.970 ;
        RECT 96.680 100.950 100.660 100.970 ;
        RECT 21.675 98.305 32.885 100.305 ;
        RECT 120.055 99.635 122.055 108.825 ;
        RECT 35.540 99.175 36.530 99.245 ;
        RECT 40.980 99.235 41.660 99.270 ;
        RECT 38.850 99.185 41.660 99.235 ;
        RECT 35.270 99.065 36.530 99.175 ;
        RECT 38.340 99.065 41.660 99.185 ;
        RECT 35.270 98.715 41.660 99.065 ;
        RECT 35.270 98.695 38.550 98.715 ;
        RECT 40.980 98.700 41.660 98.715 ;
        RECT 35.270 97.705 35.570 98.695 ;
        RECT 34.985 97.185 35.570 97.705 ;
        RECT 34.965 97.135 35.570 97.185 ;
        RECT 34.965 96.805 35.305 97.135 ;
        RECT 19.000 93.985 19.520 93.995 ;
        RECT 19.000 93.385 19.670 93.985 ;
        RECT 25.910 93.680 26.250 94.060 ;
        RECT 39.260 94.015 40.630 95.115 ;
        RECT 39.260 93.965 40.570 94.015 ;
        RECT 19.260 93.235 19.670 93.385 ;
        RECT 19.260 93.025 19.680 93.235 ;
        RECT 25.930 93.160 26.230 93.680 ;
        RECT 18.230 92.985 19.680 93.025 ;
        RECT 18.210 92.765 19.680 92.985 ;
        RECT 18.210 92.705 19.670 92.765 ;
        RECT 18.210 92.635 18.650 92.705 ;
        RECT 18.210 91.065 18.640 92.635 ;
        RECT 18.210 90.745 19.820 91.065 ;
        RECT 18.220 90.555 19.820 90.745 ;
        RECT 28.330 90.560 39.540 92.560 ;
        RECT 19.210 90.115 19.820 90.555 ;
        RECT 19.230 89.990 19.810 90.115 ;
        RECT 37.540 81.370 39.540 90.560 ;
        RECT 42.290 88.610 53.290 99.610 ;
        RECT 42.790 84.610 46.790 88.610 ;
        RECT 90.310 87.820 101.310 98.820 ;
        RECT 102.070 98.565 102.750 98.600 ;
        RECT 102.070 98.515 104.880 98.565 ;
        RECT 102.070 98.395 105.390 98.515 ;
        RECT 107.200 98.505 108.190 98.575 ;
        RECT 107.200 98.395 108.460 98.505 ;
        RECT 102.070 98.045 108.460 98.395 ;
        RECT 102.070 98.030 102.750 98.045 ;
        RECT 105.180 98.025 108.460 98.045 ;
        RECT 108.160 97.035 108.460 98.025 ;
        RECT 110.845 97.635 122.055 99.635 ;
        RECT 108.160 96.515 108.745 97.035 ;
        RECT 108.160 96.465 108.765 96.515 ;
        RECT 108.425 96.135 108.765 96.465 ;
        RECT 103.100 93.345 104.470 94.445 ;
        RECT 103.160 93.295 104.470 93.345 ;
        RECT 117.480 93.010 117.820 93.390 ;
        RECT 124.210 93.315 124.730 93.325 ;
        RECT 117.500 92.490 117.800 93.010 ;
        RECT 124.060 92.715 124.730 93.315 ;
        RECT 124.060 92.565 124.470 92.715 ;
        RECT 124.050 92.355 124.470 92.565 ;
        RECT 124.050 92.315 125.500 92.355 ;
        RECT 124.050 92.095 125.520 92.315 ;
        RECT 124.060 92.035 125.520 92.095 ;
        RECT 125.080 91.965 125.520 92.035 ;
        RECT 104.190 89.890 115.400 91.890 ;
        RECT 125.090 90.395 125.520 91.965 ;
        RECT 123.910 90.075 125.520 90.395 ;
        RECT 96.810 83.820 100.810 87.820 ;
        RECT 104.190 80.700 106.190 89.890 ;
        RECT 123.910 89.885 125.510 90.075 ;
        RECT 123.910 89.445 124.520 89.885 ;
        RECT 123.920 89.320 124.500 89.445 ;
        RECT 42.270 63.090 46.310 77.800 ;
        RECT 42.270 63.010 57.190 63.090 ;
        RECT 21.345 49.735 23.345 58.925 ;
        RECT 42.270 56.630 68.080 63.010 ;
        RECT 42.270 56.590 72.100 56.630 ;
        RECT 42.190 52.650 72.100 56.590 ;
        RECT 42.190 52.590 72.080 52.650 ;
        RECT 46.190 52.510 72.080 52.590 ;
        RECT 46.190 52.090 68.080 52.510 ;
        RECT 57.080 52.010 68.080 52.090 ;
        RECT 119.395 49.735 121.395 58.925 ;
        RECT 21.345 47.735 32.555 49.735 ;
        RECT 35.210 48.605 36.200 48.675 ;
        RECT 40.650 48.665 41.330 48.700 ;
        RECT 38.520 48.615 41.330 48.665 ;
        RECT 34.940 48.495 36.200 48.605 ;
        RECT 38.010 48.495 41.330 48.615 ;
        RECT 34.940 48.145 41.330 48.495 ;
        RECT 34.940 48.125 38.220 48.145 ;
        RECT 40.650 48.130 41.330 48.145 ;
        RECT 34.940 47.135 35.240 48.125 ;
        RECT 34.655 46.615 35.240 47.135 ;
        RECT 34.635 46.565 35.240 46.615 ;
        RECT 34.635 46.235 34.975 46.565 ;
        RECT 18.670 43.415 19.190 43.425 ;
        RECT 18.670 42.815 19.340 43.415 ;
        RECT 25.580 43.110 25.920 43.490 ;
        RECT 38.930 43.445 40.300 44.545 ;
        RECT 38.930 43.395 40.240 43.445 ;
        RECT 18.930 42.665 19.340 42.815 ;
        RECT 18.930 42.455 19.350 42.665 ;
        RECT 25.600 42.590 25.900 43.110 ;
        RECT 17.900 42.415 19.350 42.455 ;
        RECT 17.880 42.195 19.350 42.415 ;
        RECT 17.880 42.135 19.340 42.195 ;
        RECT 17.880 42.065 18.320 42.135 ;
        RECT 17.880 40.495 18.310 42.065 ;
        RECT 17.880 40.175 19.490 40.495 ;
        RECT 17.890 39.985 19.490 40.175 ;
        RECT 28.000 39.990 39.210 41.990 ;
        RECT 18.880 39.545 19.490 39.985 ;
        RECT 18.900 39.420 19.480 39.545 ;
        RECT 37.210 30.800 39.210 39.990 ;
        RECT 41.780 38.010 52.780 49.010 ;
        RECT 42.280 34.010 46.280 38.010 ;
        RECT 89.300 37.990 100.300 48.990 ;
        RECT 101.410 48.665 102.090 48.700 ;
        RECT 101.410 48.615 104.220 48.665 ;
        RECT 101.410 48.495 104.730 48.615 ;
        RECT 106.540 48.605 107.530 48.675 ;
        RECT 106.540 48.495 107.800 48.605 ;
        RECT 101.410 48.145 107.800 48.495 ;
        RECT 101.410 48.130 102.090 48.145 ;
        RECT 104.520 48.125 107.800 48.145 ;
        RECT 107.500 47.135 107.800 48.125 ;
        RECT 110.185 47.735 121.395 49.735 ;
        RECT 107.500 46.615 108.085 47.135 ;
        RECT 107.500 46.565 108.105 46.615 ;
        RECT 107.765 46.235 108.105 46.565 ;
        RECT 102.440 43.445 103.810 44.545 ;
        RECT 102.500 43.395 103.810 43.445 ;
        RECT 116.820 43.110 117.160 43.490 ;
        RECT 123.550 43.415 124.070 43.425 ;
        RECT 116.840 42.590 117.140 43.110 ;
        RECT 123.400 42.815 124.070 43.415 ;
        RECT 123.400 42.665 123.810 42.815 ;
        RECT 123.390 42.455 123.810 42.665 ;
        RECT 123.390 42.415 124.840 42.455 ;
        RECT 123.390 42.195 124.860 42.415 ;
        RECT 123.400 42.135 124.860 42.195 ;
        RECT 124.420 42.065 124.860 42.135 ;
        RECT 103.530 39.990 114.740 41.990 ;
        RECT 124.430 40.495 124.860 42.065 ;
        RECT 123.250 40.175 124.860 40.495 ;
        RECT 95.800 33.990 99.800 37.990 ;
        RECT 40.990 21.790 51.990 32.790 ;
        RECT 103.530 30.800 105.530 39.990 ;
        RECT 123.250 39.985 124.850 40.175 ;
        RECT 123.250 39.545 123.860 39.985 ;
        RECT 123.260 39.420 123.840 39.545 ;
        RECT 47.490 17.790 51.490 21.790 ;
      LAYER met4 ;
        RECT 78.850 211.400 82.860 213.760 ;
        RECT 78.850 209.660 85.570 211.400 ;
        RECT 66.540 209.580 85.570 209.660 ;
        RECT 47.640 209.500 85.570 209.580 ;
        RECT 47.640 204.580 88.430 209.500 ;
        RECT 29.425 194.695 30.325 198.105 ;
        RECT 29.425 194.605 30.330 194.695 ;
        RECT 29.480 191.860 30.330 194.605 ;
        RECT 29.480 191.725 30.470 191.860 ;
        RECT 29.570 189.865 30.470 191.725 ;
        RECT 38.660 189.865 39.500 192.905 ;
        RECT 47.640 192.330 52.640 204.580 ;
        RECT 66.540 204.500 88.430 204.580 ;
        RECT 66.540 204.460 85.570 204.500 ;
        RECT 78.850 202.730 85.570 204.460 ;
        RECT 78.850 200.530 82.860 202.730 ;
        RECT 91.195 199.495 95.325 203.625 ;
        RECT 91.200 192.370 95.320 199.495 ;
        RECT 112.745 194.695 113.645 198.105 ;
        RECT 112.740 194.605 113.645 194.695 ;
        RECT 29.570 188.995 39.500 189.865 ;
        RECT 29.570 188.360 30.470 188.995 ;
        RECT 38.660 188.945 39.500 188.995 ;
        RECT 47.240 189.010 52.640 192.330 ;
        RECT 47.240 186.390 52.240 189.010 ;
        RECT 47.180 183.965 58.540 186.390 ;
        RECT 47.180 182.270 61.255 183.965 ;
        RECT 90.850 182.370 95.850 192.370 ;
        RECT 103.570 189.865 104.410 192.905 ;
        RECT 112.740 191.860 113.590 194.605 ;
        RECT 112.600 191.725 113.590 191.860 ;
        RECT 112.600 189.865 113.500 191.725 ;
        RECT 103.570 188.995 113.500 189.865 ;
        RECT 103.570 188.945 104.410 188.995 ;
        RECT 112.600 188.360 113.500 188.995 ;
        RECT 46.780 177.310 51.780 180.170 ;
        RECT 54.420 179.840 61.255 182.270 ;
        RECT 57.125 179.835 61.255 179.840 ;
        RECT 91.210 180.910 95.315 182.370 ;
        RECT 91.210 178.050 96.290 180.910 ;
        RECT 44.880 174.600 53.550 177.310 ;
        RECT 89.390 175.340 98.060 178.050 ;
        RECT 42.520 170.590 55.750 174.600 ;
        RECT 87.030 171.330 100.260 175.340 ;
        RECT 46.620 158.280 51.820 170.590 ;
        RECT 91.130 159.020 96.330 171.330 ;
        RECT 29.425 145.125 30.325 148.535 ;
        RECT 29.425 145.035 30.330 145.125 ;
        RECT 29.480 142.290 30.330 145.035 ;
        RECT 29.480 142.155 30.470 142.290 ;
        RECT 29.570 140.295 30.470 142.155 ;
        RECT 38.660 140.295 39.500 143.335 ;
        RECT 29.570 139.425 39.500 140.295 ;
        RECT 29.570 138.790 30.470 139.425 ;
        RECT 38.660 139.375 39.500 139.425 ;
        RECT 46.700 142.800 51.700 158.280 ;
        RECT 91.210 151.020 96.210 159.020 ;
        RECT 112.745 145.125 113.645 148.535 ;
        RECT 112.740 145.035 113.645 145.125 ;
        RECT 46.700 137.010 52.290 142.800 ;
        RECT 84.265 142.110 88.315 142.115 ;
        RECT 90.720 142.110 95.720 142.760 ;
        RECT 84.265 138.070 95.720 142.110 ;
        RECT 103.570 140.295 104.410 143.335 ;
        RECT 112.740 142.290 113.590 145.035 ;
        RECT 112.600 142.155 113.590 142.290 ;
        RECT 112.600 140.295 113.500 142.155 ;
        RECT 103.570 139.425 113.500 140.295 ;
        RECT 103.570 139.375 104.410 139.425 ;
        RECT 112.600 138.790 113.500 139.425 ;
        RECT 84.265 138.065 88.315 138.070 ;
        RECT 46.700 137.000 56.250 137.010 ;
        RECT 47.290 132.800 56.250 137.000 ;
        RECT 46.250 123.830 51.250 131.830 ;
        RECT 52.210 131.755 56.250 132.800 ;
        RECT 52.205 127.705 56.255 131.755 ;
        RECT 46.170 111.520 51.370 123.830 ;
        RECT 90.720 122.860 95.720 138.070 ;
        RECT 42.070 107.510 55.300 111.520 ;
        RECT 90.640 110.550 95.840 122.860 ;
        RECT 44.430 104.800 53.100 107.510 ;
        RECT 86.540 106.540 99.770 110.550 ;
        RECT 46.330 101.940 51.710 104.800 ;
        RECT 30.085 96.895 30.985 100.305 ;
        RECT 30.085 96.805 30.990 96.895 ;
        RECT 30.140 94.060 30.990 96.805 ;
        RECT 30.140 93.925 31.130 94.060 ;
        RECT 30.230 92.065 31.130 93.925 ;
        RECT 39.320 92.065 40.160 95.105 ;
        RECT 47.770 94.610 51.710 101.940 ;
        RECT 83.455 100.965 87.585 105.095 ;
        RECT 88.900 103.830 97.570 106.540 ;
        RECT 90.800 100.970 95.800 103.830 ;
        RECT 83.460 97.520 87.580 100.965 ;
        RECT 47.770 92.340 52.790 94.610 ;
        RECT 83.460 93.400 96.020 97.520 ;
        RECT 112.745 96.225 113.645 99.635 ;
        RECT 112.740 96.135 113.645 96.225 ;
        RECT 30.230 91.195 40.160 92.065 ;
        RECT 30.230 90.560 31.130 91.195 ;
        RECT 39.320 91.145 40.160 91.195 ;
        RECT 47.790 84.610 52.790 92.340 ;
        RECT 90.810 89.140 96.020 93.400 ;
        RECT 103.570 91.395 104.410 94.435 ;
        RECT 112.740 93.390 113.590 96.135 ;
        RECT 112.600 93.255 113.590 93.390 ;
        RECT 112.600 91.395 113.500 93.255 ;
        RECT 103.570 90.525 113.500 91.395 ;
        RECT 103.570 90.475 104.410 90.525 ;
        RECT 112.600 89.890 113.500 90.525 ;
        RECT 42.265 77.770 46.315 77.775 ;
        RECT 48.730 77.770 52.770 84.610 ;
        RECT 77.010 79.150 81.020 81.510 ;
        RECT 42.265 73.730 52.770 77.770 ;
        RECT 74.300 77.410 81.020 79.150 ;
        RECT 90.810 77.410 95.810 89.140 ;
        RECT 74.300 77.330 95.810 77.410 ;
        RECT 74.300 77.250 101.330 77.330 ;
        RECT 42.265 73.725 46.315 73.730 ;
        RECT 71.440 72.330 101.330 77.250 ;
        RECT 71.440 72.250 93.330 72.330 ;
        RECT 74.300 72.210 93.330 72.250 ;
        RECT 74.300 70.480 81.020 72.210 ;
        RECT 77.010 68.280 81.020 70.480 ;
        RECT 62.500 64.410 66.510 66.770 ;
        RECT 47.080 62.670 52.130 62.750 ;
        RECT 62.500 62.670 69.220 64.410 ;
        RECT 47.080 62.590 69.220 62.670 ;
        RECT 42.190 62.510 69.220 62.590 ;
        RECT 42.190 57.590 72.080 62.510 ;
        RECT 47.080 57.510 72.080 57.590 ;
        RECT 47.080 57.470 69.220 57.510 ;
        RECT 29.755 46.325 30.655 49.735 ;
        RECT 29.755 46.235 30.660 46.325 ;
        RECT 29.810 43.490 30.660 46.235 ;
        RECT 29.810 43.355 30.800 43.490 ;
        RECT 29.900 41.495 30.800 43.355 ;
        RECT 38.990 41.495 39.830 44.535 ;
        RECT 29.900 40.625 39.830 41.495 ;
        RECT 29.900 39.990 30.800 40.625 ;
        RECT 38.990 40.575 39.830 40.625 ;
        RECT 47.080 44.010 52.130 57.470 ;
        RECT 62.500 55.740 69.220 57.470 ;
        RECT 62.500 53.540 66.510 55.740 ;
        RECT 112.085 46.325 112.985 49.735 ;
        RECT 112.080 46.235 112.985 46.325 ;
        RECT 47.080 39.800 52.280 44.010 ;
        RECT 102.910 41.495 103.750 44.535 ;
        RECT 112.080 43.490 112.930 46.235 ;
        RECT 111.940 43.355 112.930 43.490 ;
        RECT 111.940 41.495 112.840 43.355 ;
        RECT 102.910 40.625 112.840 41.495 ;
        RECT 102.910 40.575 103.750 40.625 ;
        RECT 111.940 39.990 112.840 40.625 ;
        RECT 47.280 34.010 52.280 39.800 ;
        RECT 47.390 18.320 51.450 34.010 ;
        RECT 47.390 18.220 51.270 18.320 ;
  END
END tt_um_veswaranandam_saradc_dac
END LIBRARY

