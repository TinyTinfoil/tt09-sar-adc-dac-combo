magic
tech sky130A
magscale 1 2
timestamp 1731256823
<< metal1 >>
rect 8016 38574 8584 38587
rect 8016 38372 9118 38574
rect 8348 38360 9118 38372
rect 8568 37206 8976 38360
rect 8568 36870 8614 37206
rect 8910 36870 8976 37206
rect 8568 36794 8976 36870
rect 8058 28668 8508 28675
rect 8058 28460 9128 28668
rect 8358 28454 9128 28460
rect 8578 27300 8986 28454
rect 8578 26964 8624 27300
rect 8920 26964 8986 27300
rect 8578 26888 8986 26964
rect 8314 19030 8522 19036
rect 8314 18816 9228 19030
rect 8314 18814 8522 18816
rect 8678 17662 9086 18816
rect 8678 17326 8724 17662
rect 9020 17326 9086 17662
rect 8678 17250 9086 17326
rect 4123 14069 4325 14075
rect 10913 14069 11115 43452
rect 20118 38582 20500 38586
rect 19500 38384 20500 38582
rect 19500 38368 20270 38384
rect 19642 37214 20050 38368
rect 19642 36878 19708 37214
rect 20004 36878 20050 37214
rect 19642 36802 20050 36878
rect 20034 28660 20590 28670
rect 19474 28468 20590 28660
rect 19474 28446 20244 28468
rect 19616 27292 20024 28446
rect 19616 26956 19682 27292
rect 19978 26956 20024 27292
rect 19616 26880 20024 26956
rect 19994 18872 20634 18878
rect 19492 18676 20634 18872
rect 19492 18658 20262 18676
rect 19634 17504 20042 18658
rect 19634 17168 19700 17504
rect 19996 17168 20042 17504
rect 19634 17092 20042 17168
rect 4325 13867 11115 14069
rect 4123 13861 4325 13867
rect 8188 8696 9126 8910
rect 19876 8906 20450 8938
rect 8576 7542 8984 8696
rect 19290 8692 20450 8906
rect 8576 7206 8622 7542
rect 8918 7206 8984 7542
rect 8576 7130 8984 7206
rect 19432 7538 19840 8692
rect 19876 8682 20450 8692
rect 19432 7202 19498 7538
rect 19794 7202 19840 7538
rect 19432 7126 19840 7202
rect 5116 2242 25212 2671
<< via1 >>
rect 8614 36870 8910 37206
rect 8624 26964 8920 27300
rect 8724 17326 9020 17662
rect 19708 36878 20004 37214
rect 19682 26956 19978 27292
rect 19700 17168 19996 17504
rect 4123 13867 4325 14069
rect 8622 7206 8918 7542
rect 19498 7202 19794 7538
<< metal2 >>
rect 8532 37262 9140 37288
rect 8486 37252 9186 37262
rect 8486 36594 9186 36604
rect 11388 36051 11623 43452
rect 7947 35816 11623 36051
rect 7947 33691 8182 35816
rect 12243 34997 12445 43452
rect 10775 34795 12445 34997
rect 7944 33469 7953 33691
rect 8175 33469 8184 33691
rect 7947 33463 8182 33469
rect 8542 27356 9150 27382
rect 8496 27346 9196 27356
rect 8496 26688 9196 26698
rect 3023 23937 3215 23941
rect 10775 23937 10977 34795
rect 3018 23932 10977 23937
rect 3018 23740 3023 23932
rect 3215 23740 10977 23932
rect 3018 23735 10977 23740
rect 3023 23731 3215 23735
rect 15099 21903 15301 43452
rect 20107 40991 20309 43452
rect 16621 40789 20309 40991
rect 16621 23877 16823 40789
rect 19478 37270 20086 37296
rect 19432 37260 20132 37270
rect 19432 36602 20132 36612
rect 19452 27348 20060 27374
rect 19406 27338 20106 27348
rect 19406 26680 20106 26690
rect 24752 23877 24944 23881
rect 16621 23872 24949 23877
rect 16621 23680 24752 23872
rect 24944 23680 24949 23872
rect 16621 23675 24949 23680
rect 24752 23671 24944 23675
rect 15099 21701 16713 21903
rect 8642 17718 9250 17744
rect 8596 17708 9296 17718
rect 8596 17050 9296 17060
rect 2952 14064 4123 14069
rect 2948 13872 2957 14064
rect 3149 13872 4123 14064
rect 2952 13867 4123 13872
rect 4325 13867 4331 14069
rect 16511 14047 16713 21701
rect 19470 17560 20078 17586
rect 19424 17550 20124 17560
rect 19424 16892 20124 16902
rect 16511 13845 25212 14047
rect 8540 7598 9148 7624
rect 8494 7588 9194 7598
rect 19268 7594 19876 7620
rect 8494 6930 9194 6940
rect 19222 7584 19922 7594
rect 19222 6926 19922 6936
rect 5116 2282 25212 2778
<< via2 >>
rect 8486 37206 9186 37252
rect 8486 36870 8614 37206
rect 8614 36870 8910 37206
rect 8910 36870 9186 37206
rect 8486 36604 9186 36870
rect 7953 33469 8175 33691
rect 8496 27300 9196 27346
rect 8496 26964 8624 27300
rect 8624 26964 8920 27300
rect 8920 26964 9196 27300
rect 8496 26698 9196 26964
rect 3023 23740 3215 23932
rect 19432 37214 20132 37260
rect 19432 36878 19708 37214
rect 19708 36878 20004 37214
rect 20004 36878 20132 37214
rect 19432 36612 20132 36878
rect 19406 27292 20106 27338
rect 19406 26956 19682 27292
rect 19682 26956 19978 27292
rect 19978 26956 20106 27292
rect 19406 26690 20106 26956
rect 24752 23680 24944 23872
rect 8596 17662 9296 17708
rect 8596 17326 8724 17662
rect 8724 17326 9020 17662
rect 9020 17326 9296 17662
rect 8596 17060 9296 17326
rect 2957 13872 3149 14064
rect 19424 17504 20124 17550
rect 19424 17168 19700 17504
rect 19700 17168 19996 17504
rect 19996 17168 20124 17504
rect 19424 16902 20124 17168
rect 8494 7542 9194 7588
rect 8494 7206 8622 7542
rect 8622 7206 8918 7542
rect 8918 7206 9194 7542
rect 8494 6940 9194 7206
rect 19222 7538 19922 7584
rect 19222 7202 19498 7538
rect 19498 7202 19794 7538
rect 19794 7202 19922 7538
rect 19222 6936 19922 7202
<< metal3 >>
rect 2864 43512 3042 43514
rect 2864 43452 9610 43512
rect 2864 43304 24662 43452
rect 2864 39502 3042 43304
rect 16862 39900 18240 40724
rect 19064 39900 19070 40724
rect 8348 37266 10548 39466
rect 18070 37274 20270 39474
rect 8448 37252 9248 37266
rect 8448 36604 8486 37252
rect 9186 36604 9248 37252
rect 19370 37260 20170 37274
rect 8448 36466 9248 36604
rect 10532 35968 11426 36792
rect 12250 35968 12256 36792
rect 19370 36612 19432 37260
rect 20132 36612 20170 37260
rect 19370 36474 20170 36612
rect 10532 35206 11356 35968
rect 2296 33691 8318 33696
rect 2296 33469 7953 33691
rect 8175 33469 8318 33691
rect 2296 33464 8318 33469
rect 2296 29602 2528 33464
rect 16854 30220 20242 31028
rect 8358 27360 10558 29560
rect 16854 28422 17662 30220
rect 16854 27608 17662 27614
rect 8458 27346 9258 27360
rect 18044 27352 20244 29552
rect 8458 26698 8496 27346
rect 9196 26698 9258 27346
rect 8458 26560 9258 26698
rect 19344 27338 20144 27352
rect 19344 26690 19406 27338
rect 20106 26690 20144 27338
rect 19344 26552 20144 26690
rect 10442 26350 11250 26356
rect 10442 25536 11250 25542
rect 3018 23932 3220 23937
rect 3018 23740 3023 23932
rect 3215 23740 3220 23932
rect 3018 20716 3220 23740
rect 24747 23872 25212 23877
rect 24747 23680 24752 23872
rect 24944 23680 25212 23872
rect 24747 23675 25212 23680
rect 16692 21018 17516 21024
rect 17516 20194 20160 21018
rect 16692 20188 17516 20194
rect 8458 17722 10658 19922
rect 8558 17708 9358 17722
rect 8558 17060 8596 17708
rect 9296 17060 9358 17708
rect 18062 17564 20262 19764
rect 8558 16922 9358 17060
rect 19362 17550 20162 17564
rect 19362 16902 19424 17550
rect 20124 16902 20162 17550
rect 19362 16764 20162 16902
rect 8454 15554 9262 15560
rect 2952 14064 3154 14069
rect 2952 13872 2957 14064
rect 3149 13872 3154 14064
rect 2952 11196 3154 13872
rect 8454 10518 9262 14746
rect 19266 12338 20074 14274
rect 19260 11530 19266 12338
rect 20074 11530 20080 12338
rect 17860 7598 20060 9798
rect 8484 7588 9204 7593
rect 8484 6940 8494 7588
rect 9194 6940 9204 7588
rect 8484 6935 9204 6940
rect 19160 7584 19960 7598
rect 19160 6936 19222 7584
rect 19922 6936 19960 7584
rect 19160 6798 19960 6936
rect 9536 3690 9546 4420
rect 10204 3690 10214 4420
rect 17990 4309 18930 4310
rect 17955 3371 17961 4309
rect 18959 3371 18965 4309
rect 17990 1634 18930 3371
<< via3 >>
rect 18240 39900 19064 40724
rect 11426 35968 12250 36792
rect 16854 27614 17662 28422
rect 10442 25542 11250 26350
rect 16692 20194 17516 21018
rect 8454 14746 9262 15554
rect 19266 11530 20074 12338
rect 9546 3690 10204 4420
rect 17961 3371 18959 4309
<< mimcap >>
rect 8448 38366 10448 39366
rect 8448 37466 9548 38366
rect 10348 37466 10448 38366
rect 8448 37366 10448 37466
rect 18170 38374 20170 39374
rect 18170 37474 18270 38374
rect 19070 37474 20170 38374
rect 18170 37374 20170 37474
rect 8458 28460 10458 29460
rect 8458 27560 9558 28460
rect 10358 27560 10458 28460
rect 8458 27460 10458 27560
rect 18144 28452 20144 29452
rect 18144 27552 18244 28452
rect 19044 27552 20144 28452
rect 18144 27452 20144 27552
rect 8558 18822 10558 19822
rect 8558 17922 9658 18822
rect 10458 17922 10558 18822
rect 8558 17822 10558 17922
rect 18162 18664 20162 19664
rect 18162 17764 18262 18664
rect 19062 17764 20162 18664
rect 18162 17664 20162 17764
rect 17960 8698 19960 9698
rect 17960 7798 18060 8698
rect 18860 7798 19960 8698
rect 17960 7698 19960 7798
<< mimcapcontact >>
rect 9548 37466 10348 38366
rect 18270 37474 19070 38374
rect 9558 27560 10358 28460
rect 18244 27552 19044 28452
rect 9658 17922 10458 18822
rect 18262 17764 19062 18664
rect 18060 7798 18860 8698
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 200 1000 600 44152
rect 800 1000 1200 44152
rect 1400 1000 1800 44152
rect 9528 40916 12708 41916
rect 9528 38466 10528 40916
rect 18239 40724 19065 40725
rect 18239 39900 18240 40724
rect 19064 39900 19065 40724
rect 18239 39899 19065 39900
rect 18240 38474 19064 39899
rect 9448 38366 10528 38466
rect 9448 37466 9548 38366
rect 10348 37802 10528 38366
rect 18170 38374 19170 38474
rect 10348 37466 10448 37802
rect 9448 37278 10448 37466
rect 18170 37474 18270 38374
rect 19070 37474 19170 38374
rect 9436 36793 11708 37278
rect 9436 36792 12251 36793
rect 9436 36454 11426 36792
rect 10884 35968 11426 36454
rect 12250 35968 12251 36792
rect 18170 36474 19170 37474
rect 11425 35967 12251 35968
rect 18242 35434 19063 36474
rect 9340 28560 10340 31056
rect 9340 28460 10458 28560
rect 9340 27560 9558 28460
rect 10358 27560 10458 28460
rect 18144 28452 19144 28552
rect 16853 28422 17663 28423
rect 18144 28422 18244 28452
rect 16853 27614 16854 28422
rect 17662 27614 18244 28422
rect 16853 27613 17663 27614
rect 9340 27402 10458 27560
rect 18144 27552 18244 27614
rect 19044 27552 19144 28452
rect 9340 27400 11250 27402
rect 9458 26560 11250 27400
rect 10442 26351 11250 26560
rect 10441 26350 11251 26351
rect 10441 25542 10442 26350
rect 11250 25542 11251 26350
rect 10441 25541 11251 25542
rect 18144 25300 19144 27552
rect 9554 18922 10342 21206
rect 16691 21018 17517 21019
rect 16691 20194 16692 21018
rect 17516 20194 17517 21018
rect 16691 20193 17517 20194
rect 16692 19504 17516 20193
rect 9554 18822 10558 18922
rect 9554 18468 9658 18822
rect 9558 17922 9658 18468
rect 10458 17922 10558 18822
rect 16692 18680 19204 19504
rect 9558 16922 10558 17922
rect 18162 18664 19204 18680
rect 18162 17764 18262 18664
rect 19062 17828 19204 18664
rect 19062 17764 19162 17828
rect 8453 15554 9263 15555
rect 9746 15554 10554 16922
rect 8453 14746 8454 15554
rect 9262 14746 10554 15554
rect 8453 14745 9263 14746
rect 18162 14490 19162 17764
rect 9416 7960 10426 12550
rect 19265 12338 20075 12339
rect 18026 11530 19266 12338
rect 20074 11530 20075 12338
rect 18026 8798 18834 11530
rect 19265 11529 20075 11530
rect 17960 8698 18960 8798
rect 17960 7798 18060 8698
rect 18860 7798 18960 8698
rect 9514 7078 10290 7098
rect 8222 2790 9258 5328
rect 9478 4420 10290 7078
rect 9478 3690 9546 4420
rect 10204 3690 10290 4420
rect 9478 3664 10290 3690
rect 17960 4309 18960 7798
rect 9478 3644 10254 3664
rect 17960 3371 17961 4309
rect 18959 3371 18960 4309
rect 17960 3370 18960 3371
rect 5116 2388 25212 2790
rect 8222 2266 9258 2388
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use dacswitch  dacswitch_0
timestamp 1731256823
transform 1 0 -1940 0 1 39157
box 6104 -5137 9755 4116
use dacswitch  dacswitch_1
timestamp 1731256823
transform -1 0 30554 0 1 39157
box 6104 -5137 9755 4116
use dacswitch  dacswitch_2
timestamp 1731256823
transform 1 0 -1940 0 1 29243
box 6104 -5137 9755 4116
use dacswitch  dacswitch_3
timestamp 1731256823
transform -1 0 30554 0 1 29243
box 6104 -5137 9755 4116
use dacswitch  dacswitch_4
timestamp 1731256823
transform 1 0 -1808 0 1 19597
box 6104 -5137 9755 4116
use dacswitch  dacswitch_5
timestamp 1731256823
transform -1 0 30554 0 1 19463
box 6104 -5137 9755 4116
use dacswitch  dacswitch_6
timestamp 1731256823
transform 1 0 -1874 0 1 9483
box 6104 -5137 9755 4116
use dacswitch  dacswitch_7
timestamp 1731256823
transform -1 0 30422 0 1 9483
box 6104 -5137 9755 4116
use mim400  mim400_0
timestamp 1731256823
transform 1 0 18142 0 1 30204
box -736 0 2216 5982
use mim400  mim400_1
timestamp 1731256823
transform 1 0 9150 0 -1 26366
box -736 0 2216 5982
use mim400  mim400_2
timestamp 1731256823
transform 1 0 9240 0 1 30056
box -736 0 2216 5982
use mim400  mim400_3
timestamp 1731256823
transform 0 -1 20266 -1 0 15566
box -736 0 2216 5982
use mim400  mim400_4
timestamp 1731256823
transform 1 0 18044 0 -1 26172
box -736 0 2216 5982
use mim400  mim400_5
timestamp 1731256823
transform 0 1 8438 -1 0 12618
box -736 0 2216 5982
use mim400  mim400_6
timestamp 1731256823
transform 0 1 11708 -1 0 42016
box -736 0 2216 5982
use mimcaptut200b  mimcaptut200b_0
timestamp 1731256823
transform -1 0 8456 0 1 8502
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_1
timestamp 1731256823
transform 1 0 10298 0 1 5258
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_2
timestamp 1731256823
transform -1 0 8558 0 1 18622
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_3
timestamp 1731256823
transform -1 0 8458 0 1 28260
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_4
timestamp 1731256823
transform -1 0 8448 0 1 38166
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_5
timestamp 1731256823
transform 1 0 19960 0 1 8498
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_6
timestamp 1731256823
transform 1 0 20170 0 1 38174
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_7
timestamp 1731256823
transform 1 0 20144 0 1 28252
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_8
timestamp 1731256823
transform 1 0 20162 0 1 18464
box -2100 -1700 100 1300
<< labels >>
rlabel metal4 10058 16922 10058 16922 5 top
rlabel metal3 8958 16922 8958 16922 5 bot
rlabel metal4 9958 26560 9958 26560 5 top
rlabel metal3 8858 26560 8858 26560 5 bot
rlabel metal4 9948 36466 9948 36466 5 top
rlabel metal3 8848 36466 8848 36466 5 bot
rlabel metal4 18670 36474 18670 36474 5 top
rlabel metal3 19770 36474 19770 36474 5 bot
rlabel metal4 18644 26552 18644 26552 5 top
rlabel metal3 19744 26552 19744 26552 5 bot
rlabel metal4 18662 16764 18662 16764 5 top
rlabel metal3 19762 16764 19762 16764 5 bot
rlabel metal4 18460 6798 18460 6798 5 top
rlabel metal3 19560 6798 19560 6798 5 bot
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
