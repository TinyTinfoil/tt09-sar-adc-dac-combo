VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_veswaranandam_saradc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_veswaranandam_saradc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    PORT
      LAYER met4 ;
        RECT 7.000 5.000 9.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER met1 ;
        RECT 102.715 219.465 103.725 221.200 ;
        RECT 54.565 218.455 103.725 219.465 ;
        RECT 40.080 192.870 42.920 192.935 ;
        RECT 40.080 191.860 45.590 192.870 ;
        RECT 41.740 191.800 45.590 191.860 ;
        RECT 42.840 183.970 44.880 191.800 ;
        RECT 40.290 143.340 42.540 143.375 ;
        RECT 16.090 142.260 16.590 143.340 ;
        RECT 40.290 142.300 45.640 143.340 ;
        RECT 41.790 142.270 45.640 142.300 ;
        RECT 42.890 134.440 44.930 142.270 ;
        RECT 41.570 95.150 42.610 95.180 ;
        RECT 41.570 94.080 46.140 95.150 ;
        RECT 41.570 94.070 42.610 94.080 ;
        RECT 43.390 86.250 45.430 94.080 ;
        RECT 20.615 70.345 21.625 70.375 ;
        RECT 54.565 70.345 55.575 218.455 ;
        RECT 133.040 192.935 135.235 223.055 ;
        RECT 100.590 192.910 102.500 192.930 ;
        RECT 97.500 191.920 102.500 192.910 ;
        RECT 127.000 192.025 135.235 192.935 ;
        RECT 97.500 191.840 101.350 191.920 ;
        RECT 98.210 184.010 100.250 191.840 ;
        RECT 133.040 143.425 135.235 192.025 ;
        RECT 100.170 143.300 102.950 143.350 ;
        RECT 97.370 142.340 102.950 143.300 ;
        RECT 126.640 142.455 135.235 143.425 ;
        RECT 97.370 142.230 101.220 142.340 ;
        RECT 98.080 134.400 100.120 142.230 ;
        RECT 133.040 94.525 135.235 142.455 ;
        RECT 99.970 94.360 103.170 94.390 ;
        RECT 97.460 93.380 103.170 94.360 ;
        RECT 126.640 93.555 135.235 94.525 ;
        RECT 97.460 93.290 101.310 93.380 ;
        RECT 98.170 85.460 100.210 93.290 ;
        RECT 20.615 69.335 55.575 70.345 ;
        RECT 20.615 69.305 21.625 69.335 ;
        RECT 14.170 43.575 16.865 44.610 ;
        RECT 40.940 43.480 45.630 44.550 ;
        RECT 99.380 44.530 102.250 44.690 ;
        RECT 133.040 44.625 135.235 93.555 ;
        RECT 42.880 35.650 44.920 43.480 ;
        RECT 96.450 43.460 102.250 44.530 ;
        RECT 125.980 43.655 135.235 44.625 ;
        RECT 97.160 35.630 99.200 43.460 ;
        RECT 99.380 43.410 102.250 43.460 ;
        RECT 133.040 13.355 135.235 43.655 ;
        RECT 13.220 11.210 135.235 13.355 ;
        RECT 133.040 11.185 135.235 11.210 ;
      LAYER met2 ;
        RECT 75.450 222.875 76.550 223.885 ;
        RECT 56.895 220.680 58.160 221.855 ;
        RECT 16.090 189.240 17.120 190.220 ;
        RECT 42.660 186.310 45.700 186.440 ;
        RECT 42.430 182.970 45.930 186.310 ;
        RECT 56.940 180.255 58.115 220.680 ;
        RECT 61.170 218.645 62.270 219.655 ;
        RECT 39.735 179.080 58.115 180.255 ;
        RECT 39.735 168.455 40.910 179.080 ;
        RECT 61.215 174.985 62.225 218.645 ;
        RECT 53.875 173.975 62.225 174.985 ;
        RECT 39.720 167.345 40.920 168.455 ;
        RECT 39.735 167.315 40.910 167.345 ;
        RECT 16.090 139.825 17.405 140.775 ;
        RECT 42.710 136.780 45.750 136.910 ;
        RECT 42.480 133.440 45.980 136.780 ;
        RECT 53.875 119.685 54.885 173.975 ;
        RECT 17.290 118.675 54.885 119.685 ;
        RECT 75.495 109.515 76.505 222.875 ;
        RECT 108.395 218.795 109.405 221.200 ;
        RECT 129.750 221.125 130.710 221.145 ;
        RECT 118.680 220.115 130.735 221.125 ;
        RECT 129.750 220.095 130.710 220.115 ;
        RECT 100.535 217.785 109.405 218.795 ;
        RECT 119.705 219.345 120.715 219.390 ;
        RECT 127.655 219.345 128.615 219.365 ;
        RECT 119.705 218.335 128.640 219.345 ;
        RECT 119.705 218.290 120.715 218.335 ;
        RECT 127.655 218.315 128.615 218.335 ;
        RECT 100.535 204.955 101.545 217.785 ;
        RECT 83.105 203.945 101.545 204.955 ;
        RECT 83.105 119.385 84.115 203.945 ;
        RECT 132.315 190.185 134.805 223.135 ;
        RECT 125.650 189.265 134.805 190.185 ;
        RECT 97.390 186.350 100.430 186.480 ;
        RECT 97.160 183.010 100.660 186.350 ;
        RECT 132.315 140.615 134.805 189.265 ;
        RECT 125.790 139.695 134.805 140.615 ;
        RECT 97.260 136.740 100.300 136.870 ;
        RECT 97.030 133.400 100.530 136.740 ;
        RECT 123.760 119.385 124.720 119.405 ;
        RECT 83.105 118.375 124.745 119.385 ;
        RECT 123.760 118.355 124.720 118.375 ;
        RECT 75.495 108.505 83.565 109.515 ;
        RECT 43.210 88.590 46.250 88.720 ;
        RECT 42.980 85.250 46.480 88.590 ;
        RECT 14.760 70.320 21.655 70.345 ;
        RECT 14.740 69.360 21.655 70.320 ;
        RECT 14.760 69.335 21.655 69.360 ;
        RECT 82.555 70.235 83.565 108.505 ;
        RECT 132.315 91.715 134.805 139.695 ;
        RECT 125.770 90.795 134.805 91.715 ;
        RECT 97.350 87.800 100.390 87.930 ;
        RECT 97.120 84.460 100.620 87.800 ;
        RECT 126.995 70.235 127.955 70.255 ;
        RECT 82.555 69.225 127.980 70.235 ;
        RECT 126.995 69.205 127.955 69.225 ;
        RECT 14.170 41.085 17.585 41.980 ;
        RECT 132.315 41.815 134.805 90.795 ;
        RECT 125.010 40.895 134.805 41.815 ;
        RECT 42.700 37.990 45.740 38.120 ;
        RECT 42.470 34.650 45.970 37.990 ;
        RECT 96.340 37.970 99.380 38.100 ;
        RECT 96.110 34.630 99.610 37.970 ;
        RECT 132.315 13.890 134.805 40.895 ;
        RECT 13.220 11.410 134.805 13.890 ;
        RECT 132.315 11.405 134.805 11.410 ;
      LAYER met3 ;
        RECT 75.470 223.885 76.530 223.910 ;
        RECT 75.470 222.875 79.315 223.885 ;
        RECT 75.470 222.850 76.530 222.875 ;
        RECT 56.915 221.855 58.140 221.880 ;
        RECT 56.915 221.200 100.470 221.855 ;
        RECT 56.915 220.680 112.495 221.200 ;
        RECT 56.915 220.655 58.140 220.680 ;
        RECT 61.190 219.655 62.250 219.680 ;
        RECT 113.855 219.655 114.865 221.200 ;
        RECT 119.620 220.050 120.715 221.200 ;
        RECT 61.190 218.645 114.865 219.655 ;
        RECT 119.490 219.370 120.715 220.050 ;
        RECT 61.190 218.620 62.250 218.645 ;
        RECT 119.490 218.310 120.740 219.370 ;
        RECT 119.490 218.120 120.130 218.310 ;
        RECT 122.380 217.560 123.200 221.200 ;
        RECT 129.725 220.115 133.705 221.125 ;
        RECT 16.090 216.520 123.310 217.560 ;
        RECT 62.540 210.000 73.540 210.080 ;
        RECT 62.540 203.620 84.430 210.000 ;
        RECT 58.620 203.580 95.350 203.620 ;
        RECT 58.540 199.580 95.350 203.580 ;
        RECT 62.540 199.500 95.350 199.580 ;
        RECT 62.540 199.080 84.430 199.500 ;
        RECT 73.430 199.000 84.430 199.080 ;
        RECT 41.740 186.330 52.740 197.330 ;
        RECT 90.350 186.370 101.350 197.370 ;
        RECT 127.630 188.185 128.640 219.415 ;
        RECT 42.240 182.330 46.240 186.330 ;
        RECT 52.660 179.840 61.280 183.960 ;
        RECT 96.850 182.370 100.850 186.370 ;
        RECT 97.170 180.910 101.150 180.930 ;
        RECT 52.660 176.170 56.780 179.840 ;
        RECT 97.170 176.910 101.290 180.910 ;
        RECT 16.090 167.320 41.590 168.480 ;
        RECT 46.280 165.280 57.280 176.170 ;
        RECT 90.790 166.020 101.790 176.910 ;
        RECT 132.695 170.645 133.705 220.115 ;
        RECT 46.200 165.170 57.280 165.280 ;
        RECT 90.710 165.910 101.790 166.020 ;
        RECT 127.630 169.635 133.705 170.645 ;
        RECT 46.200 154.280 57.200 165.170 ;
        RECT 90.710 155.140 101.710 165.910 ;
        RECT 84.270 155.020 101.710 155.140 ;
        RECT 52.660 150.360 56.700 154.280 ;
        RECT 52.700 150.280 56.700 150.360 ;
        RECT 84.270 151.100 101.210 155.020 ;
        RECT 41.790 136.800 52.790 147.800 ;
        RECT 84.270 138.040 88.310 151.100 ;
        RECT 97.210 151.020 101.210 151.100 ;
        RECT 42.290 132.800 46.290 136.800 ;
        RECT 90.220 136.760 101.220 147.760 ;
        RECT 127.630 138.615 128.640 169.635 ;
        RECT 96.720 132.760 100.720 136.760 ;
        RECT 52.250 131.780 56.250 131.830 ;
        RECT 52.210 127.830 56.250 131.780 ;
        RECT 96.720 130.780 100.720 130.860 ;
        RECT 45.750 116.940 56.750 127.830 ;
        RECT 96.680 126.860 100.720 130.780 ;
        RECT 45.750 116.830 56.830 116.940 ;
        RECT 45.830 105.940 56.830 116.830 ;
        RECT 90.220 115.970 101.220 126.860 ;
        RECT 123.735 118.375 128.640 119.385 ;
        RECT 90.220 115.860 101.300 115.970 ;
        RECT 52.210 101.940 56.330 105.940 ;
        RECT 83.460 105.090 87.580 105.120 ;
        RECT 90.300 105.090 101.300 115.860 ;
        RECT 83.460 104.970 101.300 105.090 ;
        RECT 52.210 101.920 56.190 101.940 ;
        RECT 83.460 100.970 100.800 104.970 ;
        RECT 83.460 100.940 87.580 100.970 ;
        RECT 96.680 100.950 100.660 100.970 ;
        RECT 42.290 88.610 53.290 99.610 ;
        RECT 42.790 84.610 46.790 88.610 ;
        RECT 90.310 87.820 101.310 98.820 ;
        RECT 127.630 89.715 128.640 118.375 ;
        RECT 96.810 83.820 100.810 87.820 ;
        RECT 14.760 39.815 15.770 70.345 ;
        RECT 42.270 63.090 46.310 77.800 ;
        RECT 86.330 77.750 97.330 77.830 ;
        RECT 75.440 71.370 97.330 77.750 ;
        RECT 71.420 71.330 101.250 71.370 ;
        RECT 71.420 67.390 101.330 71.330 ;
        RECT 71.440 67.330 101.330 67.390 ;
        RECT 71.440 67.250 100.370 67.330 ;
        RECT 75.440 66.830 100.370 67.250 ;
        RECT 75.440 66.750 86.440 66.830 ;
        RECT 42.270 63.010 57.190 63.090 ;
        RECT 42.270 56.630 68.080 63.010 ;
        RECT 96.330 61.690 100.370 66.830 ;
        RECT 96.300 57.650 100.400 61.690 ;
        RECT 42.270 56.590 72.100 56.630 ;
        RECT 42.190 52.650 72.100 56.590 ;
        RECT 42.190 52.590 72.080 52.650 ;
        RECT 46.190 52.510 72.080 52.590 ;
        RECT 46.190 52.090 68.080 52.510 ;
        RECT 57.080 52.010 68.080 52.090 ;
        RECT 41.780 38.010 52.780 49.010 ;
        RECT 42.280 34.010 46.280 38.010 ;
        RECT 89.300 37.990 100.300 48.990 ;
        RECT 126.970 39.815 127.980 70.235 ;
        RECT 95.800 33.990 99.800 37.990 ;
        RECT 40.990 21.790 51.990 32.790 ;
        RECT 47.490 17.790 51.490 21.790 ;
        RECT 89.950 21.545 94.650 21.550 ;
        RECT 89.775 16.855 94.825 21.545 ;
        RECT 89.950 8.030 94.650 16.855 ;
        RECT 89.950 3.330 136.750 8.030 ;
      LAYER met4 ;
        RECT 78.270 223.885 79.290 223.890 ;
        RECT 78.270 222.875 100.085 223.885 ;
        RECT 78.270 222.870 79.290 222.875 ;
        RECT 99.075 220.485 100.085 222.875 ;
        RECT 105.525 220.485 106.535 221.200 ;
        RECT 99.075 219.475 106.535 220.485 ;
        RECT 78.850 211.400 82.860 213.760 ;
        RECT 78.850 209.660 85.570 211.400 ;
        RECT 66.540 209.580 85.570 209.660 ;
        RECT 47.640 209.500 85.570 209.580 ;
        RECT 47.640 204.580 88.430 209.500 ;
        RECT 16.090 193.570 18.660 194.400 ;
        RECT 47.640 192.330 52.640 204.580 ;
        RECT 66.540 204.500 88.430 204.580 ;
        RECT 66.540 204.460 85.570 204.500 ;
        RECT 78.850 202.730 85.570 204.460 ;
        RECT 78.850 200.530 82.860 202.730 ;
        RECT 91.195 199.495 95.325 203.625 ;
        RECT 91.200 192.370 95.320 199.495 ;
        RECT 131.865 194.375 133.920 223.215 ;
        RECT 124.190 193.535 133.920 194.375 ;
        RECT 47.240 189.010 52.640 192.330 ;
        RECT 47.240 186.390 52.240 189.010 ;
        RECT 47.180 183.965 58.540 186.390 ;
        RECT 47.180 182.270 61.255 183.965 ;
        RECT 90.850 182.370 95.850 192.370 ;
        RECT 46.780 177.310 51.780 180.170 ;
        RECT 54.420 179.840 61.255 182.270 ;
        RECT 57.125 179.835 61.255 179.840 ;
        RECT 91.210 180.910 95.315 182.370 ;
        RECT 91.210 178.050 96.290 180.910 ;
        RECT 44.880 174.600 53.550 177.310 ;
        RECT 89.390 175.340 98.060 178.050 ;
        RECT 42.520 170.590 55.750 174.600 ;
        RECT 87.030 171.330 100.260 175.340 ;
        RECT 46.620 158.280 51.820 170.590 ;
        RECT 91.130 159.020 96.330 171.330 ;
        RECT 16.090 143.990 18.850 144.850 ;
        RECT 46.700 142.800 51.700 158.280 ;
        RECT 91.210 151.020 96.210 159.020 ;
        RECT 131.865 144.805 133.920 193.535 ;
        RECT 124.070 143.965 133.920 144.805 ;
        RECT 46.700 137.010 52.290 142.800 ;
        RECT 84.265 142.110 88.315 142.115 ;
        RECT 90.720 142.110 95.720 142.760 ;
        RECT 84.265 138.070 95.720 142.110 ;
        RECT 84.265 138.065 88.315 138.070 ;
        RECT 46.700 137.000 56.250 137.010 ;
        RECT 47.290 132.800 56.250 137.000 ;
        RECT 46.250 123.830 51.250 131.830 ;
        RECT 52.210 131.755 56.250 132.800 ;
        RECT 52.205 127.705 56.255 131.755 ;
        RECT 46.170 111.520 51.370 123.830 ;
        RECT 90.720 122.860 95.720 138.070 ;
        RECT 42.070 107.510 55.300 111.520 ;
        RECT 90.640 110.550 95.840 122.860 ;
        RECT 44.430 104.800 53.100 107.510 ;
        RECT 86.540 106.540 99.770 110.550 ;
        RECT 46.330 101.940 51.710 104.800 ;
        RECT 47.770 94.610 51.710 101.940 ;
        RECT 83.455 100.965 87.585 105.095 ;
        RECT 88.900 103.830 97.570 106.540 ;
        RECT 90.800 100.970 95.800 103.830 ;
        RECT 83.460 97.520 87.580 100.965 ;
        RECT 47.770 92.340 52.790 94.610 ;
        RECT 83.460 93.400 96.020 97.520 ;
        RECT 131.865 95.905 133.920 143.965 ;
        RECT 124.190 95.065 133.920 95.905 ;
        RECT 47.790 84.610 52.790 92.340 ;
        RECT 90.810 89.140 96.020 93.400 ;
        RECT 42.265 77.770 46.315 77.775 ;
        RECT 48.730 77.770 52.770 84.610 ;
        RECT 77.010 79.150 81.020 81.510 ;
        RECT 42.265 73.730 52.770 77.770 ;
        RECT 74.300 77.410 81.020 79.150 ;
        RECT 90.810 77.410 95.810 89.140 ;
        RECT 74.300 77.330 95.810 77.410 ;
        RECT 74.300 77.250 101.330 77.330 ;
        RECT 42.265 73.725 46.315 73.730 ;
        RECT 71.440 72.330 101.330 77.250 ;
        RECT 71.440 72.250 93.330 72.330 ;
        RECT 74.300 72.210 93.330 72.250 ;
        RECT 74.300 70.480 81.020 72.210 ;
        RECT 77.010 68.280 81.020 70.480 ;
        RECT 62.500 64.410 66.510 66.770 ;
        RECT 47.080 62.670 52.130 62.750 ;
        RECT 62.500 62.670 69.220 64.410 ;
        RECT 47.080 62.590 69.220 62.670 ;
        RECT 42.190 62.510 69.220 62.590 ;
        RECT 42.190 57.590 72.080 62.510 ;
        RECT 96.325 61.690 100.375 61.695 ;
        RECT 47.080 57.510 72.080 57.590 ;
        RECT 90.130 57.650 100.375 61.690 ;
        RECT 47.080 57.470 69.220 57.510 ;
        RECT 14.170 45.180 18.880 46.040 ;
        RECT 47.080 44.010 52.130 57.470 ;
        RECT 62.500 55.740 69.220 57.470 ;
        RECT 62.500 53.540 66.510 55.740 ;
        RECT 47.080 39.800 52.280 44.010 ;
        RECT 90.130 43.990 94.170 57.650 ;
        RECT 96.325 57.645 100.375 57.650 ;
        RECT 131.865 46.005 133.920 95.065 ;
        RECT 123.250 45.165 133.920 46.005 ;
        RECT 47.280 34.010 52.280 39.800 ;
        RECT 41.490 26.640 46.490 27.790 ;
        RECT 41.110 17.790 46.490 26.640 ;
        RECT 47.390 18.320 51.450 34.010 ;
        RECT 47.390 18.220 51.270 18.320 ;
        RECT 41.110 13.950 46.290 17.790 ;
        RECT 89.800 16.850 94.800 43.990 ;
        RECT 131.865 13.950 133.920 45.165 ;
        RECT 13.220 11.940 133.920 13.950 ;
        RECT 41.110 11.330 46.290 11.940 ;
        RECT 131.865 11.920 133.920 11.940 ;
        RECT 132.390 2.330 137.030 8.010 ;
        RECT 136.290 1.000 137.030 2.330 ;
  END
END tt_um_veswaranandam_saradc_dac
END LIBRARY

