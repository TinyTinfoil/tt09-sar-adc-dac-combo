magic
tech sky130A
magscale 1 2
timestamp 1731255746
<< checkpaint >>
rect 140 -260 3060 45412
<< metal1 >>
rect 20543 43893 20745 44240
rect 10913 43691 20745 43893
rect 8016 38574 8584 38587
rect 8016 38372 9118 38574
rect 8348 38360 9118 38372
rect 8568 37192 8976 38360
rect 8568 36884 8640 37192
rect 8884 36884 8976 37192
rect 8568 36794 8976 36884
rect 8058 28668 8508 28675
rect 3218 28452 3318 28668
rect 8058 28460 9128 28668
rect 8358 28454 9128 28460
rect 8578 27286 8986 28454
rect 8578 26978 8650 27286
rect 8894 26978 8986 27286
rect 8578 26888 8986 26978
rect 8314 19030 8522 19036
rect 8314 18816 9228 19030
rect 8314 18814 8522 18816
rect 8678 17648 9086 18816
rect 8678 17340 8750 17648
rect 8994 17340 9086 17648
rect 8678 17250 9086 17340
rect 4123 14069 4325 14075
rect 10913 14069 11115 43691
rect 26608 38587 27047 44508
rect 20118 38582 20500 38586
rect 19500 38384 20500 38582
rect 25400 38405 27047 38587
rect 19500 38368 20270 38384
rect 19642 37200 20050 38368
rect 19642 36892 19734 37200
rect 19978 36892 20050 37200
rect 19642 36802 20050 36892
rect 26608 28685 27047 38405
rect 20034 28660 20590 28670
rect 19474 28468 20590 28660
rect 25328 28491 27047 28685
rect 19474 28446 20244 28468
rect 19616 27278 20024 28446
rect 19616 26970 19708 27278
rect 19952 26970 20024 27278
rect 19616 26880 20024 26970
rect 26608 18905 27047 28491
rect 19994 18872 20634 18878
rect 19492 18676 20634 18872
rect 25328 18711 27047 18905
rect 19492 18658 20262 18676
rect 19634 17490 20042 18658
rect 19634 17182 19726 17490
rect 19970 17182 20042 17490
rect 19634 17092 20042 17182
rect 4123 14058 11115 14069
rect 4123 13878 4134 14058
rect 4314 13878 11115 14058
rect 4123 13867 11115 13878
rect 4123 13861 4325 13867
rect 2834 8715 3373 8922
rect 8188 8696 9126 8910
rect 19876 8906 20450 8938
rect 26608 8925 27047 18711
rect 8576 7528 8984 8696
rect 19290 8692 20450 8906
rect 25196 8731 27047 8925
rect 8576 7220 8648 7528
rect 8892 7220 8984 7528
rect 8576 7130 8984 7220
rect 19432 7524 19840 8692
rect 19876 8682 20450 8692
rect 19432 7216 19524 7524
rect 19768 7216 19840 7524
rect 19432 7126 19840 7216
rect 26608 2671 27047 8731
rect 2662 2242 27047 2671
rect 26608 2237 27047 2242
<< via1 >>
rect 8640 36884 8884 37192
rect 8650 26978 8894 27286
rect 8750 17340 8994 17648
rect 19734 36892 19978 37200
rect 19708 26970 19952 27278
rect 19726 17182 19970 17490
rect 4134 13878 4314 14058
rect 8648 7220 8892 7528
rect 19524 7216 19768 7524
<< metal2 >>
rect 11379 44361 11632 44371
rect 11379 44145 11397 44361
rect 11613 44145 11632 44361
rect 11379 44136 11632 44145
rect 3218 37848 3424 38044
rect 8532 37262 9140 37288
rect 8486 37236 9186 37262
rect 8486 36620 8488 37236
rect 9184 36620 9186 37236
rect 8486 36594 9186 36620
rect 11388 36051 11623 44136
rect 12234 43898 12454 43931
rect 12234 43762 12276 43898
rect 12412 43762 12454 43898
rect 12234 43729 12454 43762
rect 7947 35816 11623 36051
rect 7947 33691 8182 35816
rect 12243 34997 12445 43729
rect 10775 34795 12445 34997
rect 7944 33688 8184 33691
rect 7944 33472 7956 33688
rect 8172 33472 8184 33688
rect 7944 33469 8184 33472
rect 7947 33463 8182 33469
rect 3218 27965 3481 28155
rect 8542 27356 9150 27382
rect 8496 27330 9196 27356
rect 8496 26714 8498 27330
rect 9194 26714 9196 27330
rect 8496 26688 9196 26714
rect 10775 23937 10977 34795
rect 3458 23735 10977 23937
rect 15099 21903 15301 44508
rect 21679 43759 21881 44240
rect 25950 44225 26142 44229
rect 23736 44192 26147 44225
rect 23736 44056 25978 44192
rect 26114 44056 26147 44192
rect 23736 44023 26147 44056
rect 25950 44019 26142 44023
rect 20107 43557 21881 43759
rect 23941 43869 24143 43878
rect 25531 43869 25723 43873
rect 23941 43836 25728 43869
rect 23941 43700 23974 43836
rect 24110 43700 25559 43836
rect 25695 43700 25728 43836
rect 23941 43667 25728 43700
rect 23941 43658 24143 43667
rect 25531 43663 25723 43667
rect 20107 40991 20309 43557
rect 16621 40789 20309 40991
rect 16621 23877 16823 40789
rect 26463 38037 26961 44508
rect 25130 37853 26961 38037
rect 19478 37270 20086 37296
rect 19432 37244 20132 37270
rect 19432 36628 19434 37244
rect 20130 36628 20132 37244
rect 19432 36602 20132 36628
rect 26463 28123 26961 37853
rect 25158 27939 26961 28123
rect 19452 27348 20060 27374
rect 19406 27322 20106 27348
rect 19406 26706 19408 27322
rect 20104 26706 20106 27322
rect 19406 26680 20106 26706
rect 24752 23877 24944 23881
rect 16621 23844 24949 23877
rect 16621 23708 24780 23844
rect 24916 23708 24949 23844
rect 16621 23675 24949 23708
rect 24752 23671 24944 23675
rect 15099 21701 16713 21903
rect 8642 17718 9250 17744
rect 8596 17692 9296 17718
rect 8596 17076 8598 17692
rect 9294 17076 9296 17692
rect 8596 17050 9296 17076
rect 2952 14064 4331 14069
rect 2948 14058 4331 14064
rect 2948 14036 4134 14058
rect 2948 13900 2985 14036
rect 3121 13900 4134 14036
rect 2948 13878 4134 13900
rect 4314 13878 4331 14058
rect 2948 13872 4331 13878
rect 2952 13867 4331 13872
rect 16511 14047 16713 21701
rect 26463 18343 26961 27939
rect 25154 18159 26961 18343
rect 19470 17560 20078 17586
rect 19424 17534 20124 17560
rect 19424 16918 19426 17534
rect 20122 16918 20124 17534
rect 19424 16892 20124 16918
rect 25399 14047 25591 14051
rect 16511 14014 25596 14047
rect 16511 13878 25427 14014
rect 25563 13878 25596 14014
rect 16511 13845 25596 13878
rect 25399 13841 25591 13845
rect 2834 8217 3517 8396
rect 26463 8363 26961 18159
rect 25002 8179 26961 8363
rect 8540 7598 9148 7624
rect 8494 7572 9194 7598
rect 19268 7594 19876 7620
rect 8494 6956 8496 7572
rect 9192 6956 9194 7572
rect 8494 6930 9194 6956
rect 19222 7568 19922 7594
rect 19222 6952 19224 7568
rect 19920 6952 19922 7568
rect 19222 6926 19922 6952
rect 26463 2778 26961 8179
rect 2662 2282 26961 2778
rect 26463 2281 26961 2282
<< via2 >>
rect 11397 44145 11613 44361
rect 8488 37192 9184 37236
rect 8488 36884 8640 37192
rect 8640 36884 8884 37192
rect 8884 36884 9184 37192
rect 8488 36620 9184 36884
rect 12276 43762 12412 43898
rect 7956 33472 8172 33688
rect 8498 27286 9194 27330
rect 8498 26978 8650 27286
rect 8650 26978 8894 27286
rect 8894 26978 9194 27286
rect 8498 26714 9194 26978
rect 25978 44056 26114 44192
rect 23974 43700 24110 43836
rect 25559 43700 25695 43836
rect 19434 37200 20130 37244
rect 19434 36892 19734 37200
rect 19734 36892 19978 37200
rect 19978 36892 20130 37200
rect 19434 36628 20130 36892
rect 19408 27278 20104 27322
rect 19408 26970 19708 27278
rect 19708 26970 19952 27278
rect 19952 26970 20104 27278
rect 19408 26706 20104 26970
rect 24780 23708 24916 23844
rect 8598 17648 9294 17692
rect 8598 17340 8750 17648
rect 8750 17340 8994 17648
rect 8994 17340 9294 17648
rect 8598 17076 9294 17340
rect 2985 13900 3121 14036
rect 19426 17490 20122 17534
rect 19426 17182 19726 17490
rect 19726 17182 19970 17490
rect 19970 17182 20122 17490
rect 19426 16918 20122 17182
rect 25427 13878 25563 14014
rect 8496 7528 9192 7572
rect 8496 7220 8648 7528
rect 8648 7220 8892 7528
rect 8892 7220 9192 7528
rect 8496 6956 9192 7220
rect 19224 7524 19920 7568
rect 19224 7216 19524 7524
rect 19524 7216 19768 7524
rect 19768 7216 19920 7524
rect 19224 6952 19920 7216
<< metal3 >>
rect 11383 44371 11628 44376
rect 11383 44361 20094 44371
rect 11383 44145 11397 44361
rect 11613 44240 20094 44361
rect 11613 44145 22499 44240
rect 11383 44136 22499 44145
rect 11383 44131 11628 44136
rect 12238 43931 12450 43936
rect 22771 43931 22973 44240
rect 23924 44010 24143 44240
rect 12238 43898 22973 43931
rect 12238 43762 12276 43898
rect 12412 43762 22973 43898
rect 12238 43729 22973 43762
rect 23898 43874 24143 44010
rect 23898 43836 24148 43874
rect 12238 43724 12450 43729
rect 23898 43700 23974 43836
rect 24110 43700 24148 43836
rect 23898 43662 24148 43700
rect 23898 43624 24026 43662
rect 24476 43512 24640 44240
rect 25945 44192 26741 44225
rect 25945 44056 25978 44192
rect 26114 44056 26741 44192
rect 25945 44023 26741 44056
rect 25526 43836 25728 43883
rect 25526 43700 25559 43836
rect 25695 43700 25728 43836
rect 3218 43304 24662 43512
rect 16862 40704 19070 40724
rect 16862 39920 18260 40704
rect 19044 39920 19070 40704
rect 16862 39900 19070 39920
rect 8348 37266 10548 39466
rect 18070 37274 20270 39474
rect 25526 37637 25728 43700
rect 8448 37236 9248 37266
rect 8448 36620 8488 37236
rect 9184 36620 9248 37236
rect 19370 37244 20170 37274
rect 8448 36466 9248 36620
rect 10532 36772 12256 36792
rect 10532 35988 11446 36772
rect 12230 35988 12256 36772
rect 19370 36628 19434 37244
rect 20130 36628 20170 37244
rect 19370 36474 20170 36628
rect 10532 35968 12256 35988
rect 10532 35206 11356 35968
rect 26539 34129 26741 44023
rect 25526 33927 26741 34129
rect 3218 33688 8318 33696
rect 3218 33472 7956 33688
rect 8172 33472 8318 33688
rect 3218 33464 8318 33472
rect 16854 30220 20242 31028
rect 8358 27360 10558 29560
rect 16854 28410 17662 30220
rect 16854 27626 16866 28410
rect 17650 27626 17662 28410
rect 16854 27608 17662 27626
rect 8458 27330 9258 27360
rect 18044 27352 20244 29552
rect 25526 27723 25728 33927
rect 8458 26714 8498 27330
rect 9194 26714 9258 27330
rect 8458 26560 9258 26714
rect 19344 27322 20144 27352
rect 19344 26706 19408 27322
rect 20104 26706 20144 27322
rect 19344 26552 20144 26706
rect 10442 26338 11250 26356
rect 10442 25554 10454 26338
rect 11238 25554 11250 26338
rect 10442 25536 11250 25554
rect 24747 23844 25728 23877
rect 24747 23708 24780 23844
rect 24916 23708 25728 23844
rect 24747 23675 25728 23708
rect 16692 21018 17516 21024
rect 16692 20998 20160 21018
rect 16692 20214 16712 20998
rect 17496 20214 20160 20998
rect 16692 20194 20160 20214
rect 16692 20188 17516 20194
rect 8458 17722 10658 19922
rect 8558 17692 9358 17722
rect 8558 17076 8598 17692
rect 9294 17076 9358 17692
rect 18062 17564 20262 19764
rect 25526 17943 25728 23675
rect 8558 16922 9358 17076
rect 19362 17534 20162 17564
rect 19362 16918 19426 17534
rect 20122 16918 20162 17534
rect 19362 16764 20162 16918
rect 8454 15542 9262 15560
rect 8454 14758 8466 15542
rect 9250 14758 9262 15542
rect 2952 14036 3154 14069
rect 2952 13900 2985 14036
rect 3121 13900 3154 14036
rect 2952 7963 3154 13900
rect 8454 10518 9262 14758
rect 19266 12338 20074 14274
rect 25394 14014 25596 14047
rect 25394 13878 25427 14014
rect 25563 13878 25596 14014
rect 19260 12326 20080 12338
rect 19260 11542 19278 12326
rect 20062 11542 20080 12326
rect 19260 11530 20080 11542
rect 17860 7598 20060 9798
rect 25394 7963 25596 13878
rect 8484 7572 9204 7593
rect 8484 6956 8496 7572
rect 9192 6956 9204 7572
rect 8484 6935 9204 6956
rect 19160 7568 19960 7598
rect 19160 6952 19224 7568
rect 19920 6952 19960 7568
rect 19160 6798 19960 6952
rect 9536 4407 10214 4420
rect 9536 3703 9563 4407
rect 10187 3703 10214 4407
rect 17990 4309 18930 4310
rect 9536 3690 10214 3703
rect 17955 4272 18965 4309
rect 17955 3408 17988 4272
rect 18932 3408 18965 4272
rect 17955 3371 18965 3408
rect 17990 2204 18930 3371
<< via3 >>
rect 18260 39920 19044 40704
rect 11446 35988 12230 36772
rect 16866 27626 17650 28410
rect 10454 25554 11238 26338
rect 16712 20214 17496 20998
rect 8466 14758 9250 15542
rect 19278 11542 20062 12326
rect 9563 3703 10187 4407
rect 17988 3408 18932 4272
<< mimcap >>
rect 8448 38348 10448 39366
rect 8448 37484 9556 38348
rect 10340 37484 10448 38348
rect 8448 37366 10448 37484
rect 18170 38356 20170 39374
rect 18170 37492 18278 38356
rect 19062 37492 20170 38356
rect 18170 37374 20170 37492
rect 8458 28442 10458 29460
rect 8458 27578 9566 28442
rect 10350 27578 10458 28442
rect 8458 27460 10458 27578
rect 18144 28434 20144 29452
rect 18144 27570 18252 28434
rect 19036 27570 20144 28434
rect 18144 27452 20144 27570
rect 8558 18804 10558 19822
rect 8558 17940 9666 18804
rect 10450 17940 10558 18804
rect 8558 17822 10558 17940
rect 18162 18646 20162 19664
rect 18162 17782 18270 18646
rect 19054 17782 20162 18646
rect 18162 17664 20162 17782
rect 17960 8680 19960 9698
rect 17960 7816 18068 8680
rect 18852 7816 19960 8680
rect 17960 7698 19960 7816
<< mimcapcontact >>
rect 9556 37484 10340 38348
rect 18278 37492 19062 38356
rect 9566 27578 10350 28442
rect 18252 27570 19036 28434
rect 9666 17940 10450 18804
rect 18270 17782 19054 18646
rect 18068 7816 18852 8680
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6870 44952 6930 45152
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 15702 44952 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 200 1000 600 44152
rect 800 1000 1200 44152
rect 1400 1000 1800 44152
rect 19815 44097 20017 44508
rect 21105 44097 21307 44240
rect 19815 43895 21307 44097
rect 9528 40916 12708 41916
rect 3218 38714 3732 38880
rect 9528 38466 10528 40916
rect 18239 40704 19065 40725
rect 18239 39920 18260 40704
rect 19044 39920 19065 40704
rect 18239 39899 19065 39920
rect 18240 38474 19064 39899
rect 26373 38875 26784 44508
rect 24838 38707 26784 38875
rect 9448 38348 10528 38466
rect 9448 37484 9556 38348
rect 10340 37802 10528 38348
rect 18170 38356 19170 38474
rect 10340 37484 10448 37802
rect 9448 37278 10448 37484
rect 18170 37492 18278 38356
rect 19062 37492 19170 38356
rect 9436 36793 11708 37278
rect 9436 36772 12251 36793
rect 9436 36454 11446 36772
rect 10884 35988 11446 36454
rect 12230 35988 12251 36772
rect 18170 36474 19170 37492
rect 10884 35968 12251 35988
rect 11425 35967 12251 35968
rect 18242 35434 19063 36474
rect 3218 28798 3770 28970
rect 9340 28560 10340 31056
rect 26373 28961 26784 38707
rect 24814 28793 26784 28961
rect 9340 28442 10458 28560
rect 9340 27578 9566 28442
rect 10350 27578 10458 28442
rect 18144 28434 19144 28552
rect 16853 28422 17663 28423
rect 18144 28422 18252 28434
rect 16853 28410 18252 28422
rect 16853 27626 16866 28410
rect 17650 27626 18252 28410
rect 16853 27614 18252 27626
rect 16853 27613 17663 27614
rect 9340 27402 10458 27578
rect 18144 27570 18252 27614
rect 19036 27570 19144 28434
rect 9340 27400 11250 27402
rect 9458 26560 11250 27400
rect 10442 26351 11250 26560
rect 10441 26338 11251 26351
rect 10441 25554 10454 26338
rect 11238 25554 11251 26338
rect 10441 25541 11251 25554
rect 18144 25300 19144 27570
rect 9554 18922 10342 21206
rect 16691 20998 17517 21019
rect 16691 20214 16712 20998
rect 17496 20214 17517 20998
rect 16691 20193 17517 20214
rect 16692 19504 17516 20193
rect 9554 18804 10558 18922
rect 9554 18468 9666 18804
rect 9558 17940 9666 18468
rect 10450 17940 10558 18804
rect 16692 18680 19204 19504
rect 26373 19181 26784 28793
rect 24838 19013 26784 19181
rect 9558 16922 10558 17940
rect 18162 18646 19204 18680
rect 18162 17782 18270 18646
rect 19054 17828 19204 18646
rect 19054 17782 19162 17828
rect 8453 15554 9263 15555
rect 9746 15554 10554 16922
rect 8453 15542 10554 15554
rect 8453 14758 8466 15542
rect 9250 14758 10554 15542
rect 8453 14746 10554 14758
rect 8453 14745 9263 14746
rect 18162 14490 19162 17782
rect 2834 9036 3776 9208
rect 9416 7960 10426 12550
rect 19265 12338 20075 12339
rect 18026 12326 20075 12338
rect 18026 11542 19278 12326
rect 20062 11542 20075 12326
rect 18026 11530 20075 11542
rect 18026 8798 18834 11530
rect 19265 11529 20075 11530
rect 26373 9201 26784 19013
rect 24650 9033 26784 9201
rect 17960 8680 18960 8798
rect 17960 7816 18068 8680
rect 18852 7816 18960 8680
rect 9514 7078 10290 7098
rect 8222 2790 9258 5328
rect 9478 4407 10290 7078
rect 9478 3703 9563 4407
rect 10187 3703 10290 4407
rect 9478 3664 10290 3703
rect 17960 4272 18960 7816
rect 9478 3644 10254 3664
rect 17960 3408 17988 4272
rect 18932 3408 18960 4272
rect 17960 3370 18960 3408
rect 26373 2790 26784 9033
rect 2662 2388 26784 2790
rect 8222 2266 9258 2388
rect 26373 2384 26784 2388
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 200
use mim400  mim400_0
timestamp 1559856578
transform 1 0 18142 0 1 30204
box -736 0 2216 5982
use mim400  mim400_1
timestamp 1559856578
transform 1 0 9150 0 -1 26366
box -736 0 2216 5982
use mim400  mim400_2
timestamp 1559856578
transform 1 0 9240 0 1 30056
box -736 0 2216 5982
use mim400  mim400_3
timestamp 1559856578
transform 0 -1 20266 -1 0 15566
box -736 0 2216 5982
use mim400  mim400_4
timestamp 1559856578
transform 1 0 18044 0 -1 26172
box -736 0 2216 5982
use mim400  mim400_5
timestamp 1559856578
transform 0 1 8438 -1 0 12618
box -736 0 2216 5982
use mim400  mim400_6
timestamp 1559856578
transform 0 1 11708 -1 0 42016
box -736 0 2216 5982
use mimcaptut200b  mimcaptut200b_0
timestamp 1559856578
transform -1 0 8456 0 1 8502
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_1
timestamp 1559856578
transform 1 0 10298 0 1 5258
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_2
timestamp 1559856578
transform -1 0 8558 0 1 18622
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_3
timestamp 1559856578
transform -1 0 8458 0 1 28260
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_4
timestamp 1559856578
transform -1 0 8448 0 1 38166
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_5
timestamp 1559856578
transform 1 0 19960 0 1 8498
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_6
timestamp 1559856578
transform 1 0 20170 0 1 38174
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_7
timestamp 1559856578
transform 1 0 20144 0 1 28252
box -2100 -1700 100 1300
use mimcaptut200b  mimcaptut200b_8
timestamp 1559856578
transform 1 0 20162 0 1 18464
box -2100 -1700 100 1300
<< labels >>
rlabel metal4 s 10058 16922 10058 16922 4 top
rlabel metal4 s 9958 26560 9958 26560 4 top
rlabel metal4 s 9948 36466 9948 36466 4 top
rlabel metal4 s 18670 36474 18670 36474 4 top
rlabel metal4 s 18644 26552 18644 26552 4 top
rlabel metal4 s 18662 16764 18662 16764 4 top
rlabel metal4 s 18460 6798 18460 6798 4 top
rlabel metal3 s 8958 16922 8958 16922 4 bot
rlabel metal3 s 8858 26560 8858 26560 4 bot
rlabel metal3 s 8848 36466 8848 36466 4 bot
rlabel metal3 s 19770 36474 19770 36474 4 bot
rlabel metal3 s 19744 26552 19744 26552 4 bot
rlabel metal3 s 19762 16764 19762 16764 4 bot
rlabel metal3 s 19560 6798 19560 6798 4 bot
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
